// nios_fprint.v

// Generated using ACDS version 13.1 162 at 2015.09.11.16:57:50

`timescale 1 ps / 1 ps
module nios_fprint (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire         cfpu_0_irq_export;                                                  // cfpu_0:irq -> processorM_0:fprint_irq_0_irq_export
	wire         mm_interconnect_0_memory_0_mm_bridge_0_s0_waitrequest;              // memory_0:mm_bridge_0_s0_waitrequest -> mm_interconnect_0:memory_0_mm_bridge_0_s0_waitrequest
	wire   [0:0] mm_interconnect_0_memory_0_mm_bridge_0_s0_burstcount;               // mm_interconnect_0:memory_0_mm_bridge_0_s0_burstcount -> memory_0:mm_bridge_0_s0_burstcount
	wire  [31:0] mm_interconnect_0_memory_0_mm_bridge_0_s0_writedata;                // mm_interconnect_0:memory_0_mm_bridge_0_s0_writedata -> memory_0:mm_bridge_0_s0_writedata
	wire  [22:0] mm_interconnect_0_memory_0_mm_bridge_0_s0_address;                  // mm_interconnect_0:memory_0_mm_bridge_0_s0_address -> memory_0:mm_bridge_0_s0_address
	wire         mm_interconnect_0_memory_0_mm_bridge_0_s0_write;                    // mm_interconnect_0:memory_0_mm_bridge_0_s0_write -> memory_0:mm_bridge_0_s0_write
	wire         mm_interconnect_0_memory_0_mm_bridge_0_s0_read;                     // mm_interconnect_0:memory_0_mm_bridge_0_s0_read -> memory_0:mm_bridge_0_s0_read
	wire  [31:0] mm_interconnect_0_memory_0_mm_bridge_0_s0_readdata;                 // memory_0:mm_bridge_0_s0_readdata -> mm_interconnect_0:memory_0_mm_bridge_0_s0_readdata
	wire         mm_interconnect_0_memory_0_mm_bridge_0_s0_debugaccess;              // mm_interconnect_0:memory_0_mm_bridge_0_s0_debugaccess -> memory_0:mm_bridge_0_s0_debugaccess
	wire         mm_interconnect_0_memory_0_mm_bridge_0_s0_readdatavalid;            // memory_0:mm_bridge_0_s0_readdatavalid -> mm_interconnect_0:memory_0_mm_bridge_0_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_memory_0_mm_bridge_0_s0_byteenable;               // mm_interconnect_0:memory_0_mm_bridge_0_s0_byteenable -> memory_0:mm_bridge_0_s0_byteenable
	wire   [0:0] mm_bridge_0_m0_burstcount;                                          // mm_bridge_0:m0_burstcount -> mm_interconnect_0:mm_bridge_0_m0_burstcount
	wire         mm_bridge_0_m0_waitrequest;                                         // mm_interconnect_0:mm_bridge_0_m0_waitrequest -> mm_bridge_0:m0_waitrequest
	wire  [24:0] mm_bridge_0_m0_address;                                             // mm_bridge_0:m0_address -> mm_interconnect_0:mm_bridge_0_m0_address
	wire  [31:0] mm_bridge_0_m0_writedata;                                           // mm_bridge_0:m0_writedata -> mm_interconnect_0:mm_bridge_0_m0_writedata
	wire         mm_bridge_0_m0_write;                                               // mm_bridge_0:m0_write -> mm_interconnect_0:mm_bridge_0_m0_write
	wire         mm_bridge_0_m0_read;                                                // mm_bridge_0:m0_read -> mm_interconnect_0:mm_bridge_0_m0_read
	wire  [31:0] mm_bridge_0_m0_readdata;                                            // mm_interconnect_0:mm_bridge_0_m0_readdata -> mm_bridge_0:m0_readdata
	wire         mm_bridge_0_m0_debugaccess;                                         // mm_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_bridge_0_m0_debugaccess
	wire   [3:0] mm_bridge_0_m0_byteenable;                                          // mm_bridge_0:m0_byteenable -> mm_interconnect_0:mm_bridge_0_m0_byteenable
	wire         mm_bridge_0_m0_readdatavalid;                                       // mm_interconnect_0:mm_bridge_0_m0_readdatavalid -> mm_bridge_0:m0_readdatavalid
	wire         mm_interconnect_0_cfpu_0_fprint_waitrequest;                        // cfpu_0:fprint_waitrequest -> mm_interconnect_0:cfpu_0_fprint_waitrequest
	wire  [31:0] mm_interconnect_0_cfpu_0_fprint_writedata;                          // mm_interconnect_0:cfpu_0_fprint_writedata -> cfpu_0:fprint_writedata
	wire   [9:0] mm_interconnect_0_cfpu_0_fprint_address;                            // mm_interconnect_0:cfpu_0_fprint_address -> cfpu_0:fprint_address
	wire         mm_interconnect_0_cfpu_0_fprint_write;                              // mm_interconnect_0:cfpu_0_fprint_write -> cfpu_0:fprint_write
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;                     // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;                    // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire         processor2_0_fingerprint_0_avalon_master_waitrequest;               // mm_interconnect_1:processor2_0_fingerprint_0_avalon_master_waitrequest -> processor2_0:fingerprint_0_avalon_master_waitrequest
	wire  [26:0] processor2_0_fingerprint_0_avalon_master_address;                   // processor2_0:fingerprint_0_avalon_master_address -> mm_interconnect_1:processor2_0_fingerprint_0_avalon_master_address
	wire  [31:0] processor2_0_fingerprint_0_avalon_master_writedata;                 // processor2_0:fingerprint_0_avalon_master_writedata -> mm_interconnect_1:processor2_0_fingerprint_0_avalon_master_writedata
	wire         processor2_0_fingerprint_0_avalon_master_write;                     // processor2_0:fingerprint_0_avalon_master_write -> mm_interconnect_1:processor2_0_fingerprint_0_avalon_master_write
	wire         processor2_0_fingerprint_0_avalon_master_read;                      // processor2_0:fingerprint_0_avalon_master_read -> mm_interconnect_1:processor2_0_fingerprint_0_avalon_master_read
	wire  [31:0] processor2_0_fingerprint_0_avalon_master_readdata;                  // mm_interconnect_1:processor2_0_fingerprint_0_avalon_master_readdata -> processor2_0:fingerprint_0_avalon_master_readdata
	wire  [27:0] mm_interconnect_1_processor5_0_dma_0_control_port_slave_writedata;  // mm_interconnect_1:processor5_0_dma_0_control_port_slave_writedata -> processor5_0:dma_0_control_port_slave_writedata
	wire   [2:0] mm_interconnect_1_processor5_0_dma_0_control_port_slave_address;    // mm_interconnect_1:processor5_0_dma_0_control_port_slave_address -> processor5_0:dma_0_control_port_slave_address
	wire         mm_interconnect_1_processor5_0_dma_0_control_port_slave_chipselect; // mm_interconnect_1:processor5_0_dma_0_control_port_slave_chipselect -> processor5_0:dma_0_control_port_slave_chipselect
	wire         mm_interconnect_1_processor5_0_dma_0_control_port_slave_write;      // mm_interconnect_1:processor5_0_dma_0_control_port_slave_write -> processor5_0:dma_0_control_port_slave_write_n
	wire  [27:0] mm_interconnect_1_processor5_0_dma_0_control_port_slave_readdata;   // processor5_0:dma_0_control_port_slave_readdata -> mm_interconnect_1:processor5_0_dma_0_control_port_slave_readdata
	wire   [0:0] processor2_0_out_system_bridge_m0_burstcount;                       // processor2_0:out_system_bridge_m0_burstcount -> mm_interconnect_1:processor2_0_out_system_bridge_m0_burstcount
	wire         processor2_0_out_system_bridge_m0_waitrequest;                      // mm_interconnect_1:processor2_0_out_system_bridge_m0_waitrequest -> processor2_0:out_system_bridge_m0_waitrequest
	wire  [26:0] processor2_0_out_system_bridge_m0_address;                          // processor2_0:out_system_bridge_m0_address -> mm_interconnect_1:processor2_0_out_system_bridge_m0_address
	wire  [31:0] processor2_0_out_system_bridge_m0_writedata;                        // processor2_0:out_system_bridge_m0_writedata -> mm_interconnect_1:processor2_0_out_system_bridge_m0_writedata
	wire         processor2_0_out_system_bridge_m0_write;                            // processor2_0:out_system_bridge_m0_write -> mm_interconnect_1:processor2_0_out_system_bridge_m0_write
	wire         processor2_0_out_system_bridge_m0_read;                             // processor2_0:out_system_bridge_m0_read -> mm_interconnect_1:processor2_0_out_system_bridge_m0_read
	wire  [31:0] processor2_0_out_system_bridge_m0_readdata;                         // mm_interconnect_1:processor2_0_out_system_bridge_m0_readdata -> processor2_0:out_system_bridge_m0_readdata
	wire         processor2_0_out_system_bridge_m0_debugaccess;                      // processor2_0:out_system_bridge_m0_debugaccess -> mm_interconnect_1:processor2_0_out_system_bridge_m0_debugaccess
	wire   [3:0] processor2_0_out_system_bridge_m0_byteenable;                       // processor2_0:out_system_bridge_m0_byteenable -> mm_interconnect_1:processor2_0_out_system_bridge_m0_byteenable
	wire         processor2_0_out_system_bridge_m0_readdatavalid;                    // mm_interconnect_1:processor2_0_out_system_bridge_m0_readdatavalid -> processor2_0:out_system_bridge_m0_readdatavalid
	wire   [0:0] processor6_0_out_system_bridge_m0_burstcount;                       // processor6_0:out_system_bridge_m0_burstcount -> mm_interconnect_1:processor6_0_out_system_bridge_m0_burstcount
	wire         processor6_0_out_system_bridge_m0_waitrequest;                      // mm_interconnect_1:processor6_0_out_system_bridge_m0_waitrequest -> processor6_0:out_system_bridge_m0_waitrequest
	wire  [26:0] processor6_0_out_system_bridge_m0_address;                          // processor6_0:out_system_bridge_m0_address -> mm_interconnect_1:processor6_0_out_system_bridge_m0_address
	wire  [31:0] processor6_0_out_system_bridge_m0_writedata;                        // processor6_0:out_system_bridge_m0_writedata -> mm_interconnect_1:processor6_0_out_system_bridge_m0_writedata
	wire         processor6_0_out_system_bridge_m0_write;                            // processor6_0:out_system_bridge_m0_write -> mm_interconnect_1:processor6_0_out_system_bridge_m0_write
	wire         processor6_0_out_system_bridge_m0_read;                             // processor6_0:out_system_bridge_m0_read -> mm_interconnect_1:processor6_0_out_system_bridge_m0_read
	wire  [31:0] processor6_0_out_system_bridge_m0_readdata;                         // mm_interconnect_1:processor6_0_out_system_bridge_m0_readdata -> processor6_0:out_system_bridge_m0_readdata
	wire         processor6_0_out_system_bridge_m0_debugaccess;                      // processor6_0:out_system_bridge_m0_debugaccess -> mm_interconnect_1:processor6_0_out_system_bridge_m0_debugaccess
	wire   [3:0] processor6_0_out_system_bridge_m0_byteenable;                       // processor6_0:out_system_bridge_m0_byteenable -> mm_interconnect_1:processor6_0_out_system_bridge_m0_byteenable
	wire         processor6_0_out_system_bridge_m0_readdatavalid;                    // mm_interconnect_1:processor6_0_out_system_bridge_m0_readdatavalid -> processor6_0:out_system_bridge_m0_readdatavalid
	wire  [31:0] mm_interconnect_1_processor4_0_cpu_irq_0_s0_writedata;              // mm_interconnect_1:processor4_0_cpu_irq_0_s0_writedata -> processor4_0:cpu_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processor4_0_cpu_irq_0_s0_address;                // mm_interconnect_1:processor4_0_cpu_irq_0_s0_address -> processor4_0:cpu_irq_0_s0_address
	wire         mm_interconnect_1_processor4_0_cpu_irq_0_s0_write;                  // mm_interconnect_1:processor4_0_cpu_irq_0_s0_write -> processor4_0:cpu_irq_0_s0_write
	wire  [31:0] mm_interconnect_1_processor2_0_cpu_irq_0_s0_writedata;              // mm_interconnect_1:processor2_0_cpu_irq_0_s0_writedata -> processor2_0:cpu_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processor2_0_cpu_irq_0_s0_address;                // mm_interconnect_1:processor2_0_cpu_irq_0_s0_address -> processor2_0:cpu_irq_0_s0_address
	wire         mm_interconnect_1_processor2_0_cpu_irq_0_s0_write;                  // mm_interconnect_1:processor2_0_cpu_irq_0_s0_write -> processor2_0:cpu_irq_0_s0_write
	wire  [27:0] mm_interconnect_1_processor2_0_dma_0_control_port_slave_writedata;  // mm_interconnect_1:processor2_0_dma_0_control_port_slave_writedata -> processor2_0:dma_0_control_port_slave_writedata
	wire   [2:0] mm_interconnect_1_processor2_0_dma_0_control_port_slave_address;    // mm_interconnect_1:processor2_0_dma_0_control_port_slave_address -> processor2_0:dma_0_control_port_slave_address
	wire         mm_interconnect_1_processor2_0_dma_0_control_port_slave_chipselect; // mm_interconnect_1:processor2_0_dma_0_control_port_slave_chipselect -> processor2_0:dma_0_control_port_slave_chipselect
	wire         mm_interconnect_1_processor2_0_dma_0_control_port_slave_write;      // mm_interconnect_1:processor2_0_dma_0_control_port_slave_write -> processor2_0:dma_0_control_port_slave_write_n
	wire  [27:0] mm_interconnect_1_processor2_0_dma_0_control_port_slave_readdata;   // processor2_0:dma_0_control_port_slave_readdata -> mm_interconnect_1:processor2_0_dma_0_control_port_slave_readdata
	wire  [31:0] mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_writedata; // mm_interconnect_1:processor2_0_cpu_oflow_irq_0_avs_oflow_writedata -> processor2_0:cpu_oflow_irq_0_avs_oflow_writedata
	wire   [7:0] mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_address;   // mm_interconnect_1:processor2_0_cpu_oflow_irq_0_avs_oflow_address -> processor2_0:cpu_oflow_irq_0_avs_oflow_address
	wire         mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_write;     // mm_interconnect_1:processor2_0_cpu_oflow_irq_0_avs_oflow_write -> processor2_0:cpu_oflow_irq_0_avs_oflow_write
	wire         mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_read;      // mm_interconnect_1:processor2_0_cpu_oflow_irq_0_avs_oflow_read -> processor2_0:cpu_oflow_irq_0_avs_oflow_read
	wire  [31:0] mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_readdata;  // processor2_0:cpu_oflow_irq_0_avs_oflow_readdata -> mm_interconnect_1:processor2_0_cpu_oflow_irq_0_avs_oflow_readdata
	wire         processor3_0_fingerprint_0_avalon_master_waitrequest;               // mm_interconnect_1:processor3_0_fingerprint_0_avalon_master_waitrequest -> processor3_0:fingerprint_0_avalon_master_waitrequest
	wire  [26:0] processor3_0_fingerprint_0_avalon_master_address;                   // processor3_0:fingerprint_0_avalon_master_address -> mm_interconnect_1:processor3_0_fingerprint_0_avalon_master_address
	wire  [31:0] processor3_0_fingerprint_0_avalon_master_writedata;                 // processor3_0:fingerprint_0_avalon_master_writedata -> mm_interconnect_1:processor3_0_fingerprint_0_avalon_master_writedata
	wire         processor3_0_fingerprint_0_avalon_master_write;                     // processor3_0:fingerprint_0_avalon_master_write -> mm_interconnect_1:processor3_0_fingerprint_0_avalon_master_write
	wire         processor3_0_fingerprint_0_avalon_master_read;                      // processor3_0:fingerprint_0_avalon_master_read -> mm_interconnect_1:processor3_0_fingerprint_0_avalon_master_read
	wire  [31:0] processor3_0_fingerprint_0_avalon_master_readdata;                  // mm_interconnect_1:processor3_0_fingerprint_0_avalon_master_readdata -> processor3_0:fingerprint_0_avalon_master_readdata
	wire         mm_interconnect_1_mm_bridge_0_s0_waitrequest;                       // mm_bridge_0:s0_waitrequest -> mm_interconnect_1:mm_bridge_0_s0_waitrequest
	wire   [0:0] mm_interconnect_1_mm_bridge_0_s0_burstcount;                        // mm_interconnect_1:mm_bridge_0_s0_burstcount -> mm_bridge_0:s0_burstcount
	wire  [31:0] mm_interconnect_1_mm_bridge_0_s0_writedata;                         // mm_interconnect_1:mm_bridge_0_s0_writedata -> mm_bridge_0:s0_writedata
	wire  [24:0] mm_interconnect_1_mm_bridge_0_s0_address;                           // mm_interconnect_1:mm_bridge_0_s0_address -> mm_bridge_0:s0_address
	wire         mm_interconnect_1_mm_bridge_0_s0_write;                             // mm_interconnect_1:mm_bridge_0_s0_write -> mm_bridge_0:s0_write
	wire         mm_interconnect_1_mm_bridge_0_s0_read;                              // mm_interconnect_1:mm_bridge_0_s0_read -> mm_bridge_0:s0_read
	wire  [31:0] mm_interconnect_1_mm_bridge_0_s0_readdata;                          // mm_bridge_0:s0_readdata -> mm_interconnect_1:mm_bridge_0_s0_readdata
	wire         mm_interconnect_1_mm_bridge_0_s0_debugaccess;                       // mm_interconnect_1:mm_bridge_0_s0_debugaccess -> mm_bridge_0:s0_debugaccess
	wire         mm_interconnect_1_mm_bridge_0_s0_readdatavalid;                     // mm_bridge_0:s0_readdatavalid -> mm_interconnect_1:mm_bridge_0_s0_readdatavalid
	wire   [3:0] mm_interconnect_1_mm_bridge_0_s0_byteenable;                        // mm_interconnect_1:mm_bridge_0_s0_byteenable -> mm_bridge_0:s0_byteenable
	wire         mm_interconnect_1_cfpu_0_csr_waitrequest;                           // cfpu_0:csr_waitrequest -> mm_interconnect_1:cfpu_0_csr_waitrequest
	wire  [31:0] mm_interconnect_1_cfpu_0_csr_writedata;                             // mm_interconnect_1:cfpu_0_csr_writedata -> cfpu_0:csr_writedata
	wire   [9:0] mm_interconnect_1_cfpu_0_csr_address;                               // mm_interconnect_1:cfpu_0_csr_address -> cfpu_0:csr_address
	wire         mm_interconnect_1_cfpu_0_csr_write;                                 // mm_interconnect_1:cfpu_0_csr_write -> cfpu_0:csr_write
	wire         mm_interconnect_1_cfpu_0_csr_read;                                  // mm_interconnect_1:cfpu_0_csr_read -> cfpu_0:csr_read
	wire  [31:0] mm_interconnect_1_cfpu_0_csr_readdata;                              // cfpu_0:csr_readdata -> mm_interconnect_1:cfpu_0_csr_readdata
	wire  [31:0] mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_writedata; // mm_interconnect_1:processor6_0_cpu_oflow_irq_0_avs_oflow_writedata -> processor6_0:cpu_oflow_irq_0_avs_oflow_writedata
	wire   [7:0] mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_address;   // mm_interconnect_1:processor6_0_cpu_oflow_irq_0_avs_oflow_address -> processor6_0:cpu_oflow_irq_0_avs_oflow_address
	wire         mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_write;     // mm_interconnect_1:processor6_0_cpu_oflow_irq_0_avs_oflow_write -> processor6_0:cpu_oflow_irq_0_avs_oflow_write
	wire         mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_read;      // mm_interconnect_1:processor6_0_cpu_oflow_irq_0_avs_oflow_read -> processor6_0:cpu_oflow_irq_0_avs_oflow_read
	wire  [31:0] mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_readdata;  // processor6_0:cpu_oflow_irq_0_avs_oflow_readdata -> mm_interconnect_1:processor6_0_cpu_oflow_irq_0_avs_oflow_readdata
	wire  [27:0] mm_interconnect_1_processor6_0_dma_0_control_port_slave_writedata;  // mm_interconnect_1:processor6_0_dma_0_control_port_slave_writedata -> processor6_0:dma_0_control_port_slave_writedata
	wire   [2:0] mm_interconnect_1_processor6_0_dma_0_control_port_slave_address;    // mm_interconnect_1:processor6_0_dma_0_control_port_slave_address -> processor6_0:dma_0_control_port_slave_address
	wire         mm_interconnect_1_processor6_0_dma_0_control_port_slave_chipselect; // mm_interconnect_1:processor6_0_dma_0_control_port_slave_chipselect -> processor6_0:dma_0_control_port_slave_chipselect
	wire         mm_interconnect_1_processor6_0_dma_0_control_port_slave_write;      // mm_interconnect_1:processor6_0_dma_0_control_port_slave_write -> processor6_0:dma_0_control_port_slave_write_n
	wire  [27:0] mm_interconnect_1_processor6_0_dma_0_control_port_slave_readdata;   // processor6_0:dma_0_control_port_slave_readdata -> mm_interconnect_1:processor6_0_dma_0_control_port_slave_readdata
	wire   [0:0] processor0_0_out_system_bridge_m0_burstcount;                       // processor0_0:out_system_bridge_m0_burstcount -> mm_interconnect_1:processor0_0_out_system_bridge_m0_burstcount
	wire         processor0_0_out_system_bridge_m0_waitrequest;                      // mm_interconnect_1:processor0_0_out_system_bridge_m0_waitrequest -> processor0_0:out_system_bridge_m0_waitrequest
	wire  [26:0] processor0_0_out_system_bridge_m0_address;                          // processor0_0:out_system_bridge_m0_address -> mm_interconnect_1:processor0_0_out_system_bridge_m0_address
	wire  [31:0] processor0_0_out_system_bridge_m0_writedata;                        // processor0_0:out_system_bridge_m0_writedata -> mm_interconnect_1:processor0_0_out_system_bridge_m0_writedata
	wire         processor0_0_out_system_bridge_m0_write;                            // processor0_0:out_system_bridge_m0_write -> mm_interconnect_1:processor0_0_out_system_bridge_m0_write
	wire         processor0_0_out_system_bridge_m0_read;                             // processor0_0:out_system_bridge_m0_read -> mm_interconnect_1:processor0_0_out_system_bridge_m0_read
	wire  [31:0] processor0_0_out_system_bridge_m0_readdata;                         // mm_interconnect_1:processor0_0_out_system_bridge_m0_readdata -> processor0_0:out_system_bridge_m0_readdata
	wire         processor0_0_out_system_bridge_m0_debugaccess;                      // processor0_0:out_system_bridge_m0_debugaccess -> mm_interconnect_1:processor0_0_out_system_bridge_m0_debugaccess
	wire   [3:0] processor0_0_out_system_bridge_m0_byteenable;                       // processor0_0:out_system_bridge_m0_byteenable -> mm_interconnect_1:processor0_0_out_system_bridge_m0_byteenable
	wire         processor0_0_out_system_bridge_m0_readdatavalid;                    // mm_interconnect_1:processor0_0_out_system_bridge_m0_readdatavalid -> processor0_0:out_system_bridge_m0_readdatavalid
	wire  [31:0] mm_interconnect_1_processor5_0_cpu_irq_0_s0_writedata;              // mm_interconnect_1:processor5_0_cpu_irq_0_s0_writedata -> processor5_0:cpu_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processor5_0_cpu_irq_0_s0_address;                // mm_interconnect_1:processor5_0_cpu_irq_0_s0_address -> processor5_0:cpu_irq_0_s0_address
	wire         mm_interconnect_1_processor5_0_cpu_irq_0_s0_write;                  // mm_interconnect_1:processor5_0_cpu_irq_0_s0_write -> processor5_0:cpu_irq_0_s0_write
	wire  [31:0] mm_interconnect_1_processor1_0_cpu1_irq_0_s0_writedata;             // mm_interconnect_1:processor1_0_cpu1_irq_0_s0_writedata -> processor1_0:cpu1_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processor1_0_cpu1_irq_0_s0_address;               // mm_interconnect_1:processor1_0_cpu1_irq_0_s0_address -> processor1_0:cpu1_irq_0_s0_address
	wire         mm_interconnect_1_processor1_0_cpu1_irq_0_s0_write;                 // mm_interconnect_1:processor1_0_cpu1_irq_0_s0_write -> processor1_0:cpu1_irq_0_s0_write
	wire  [31:0] mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_writedata; // mm_interconnect_1:processor7_0_cpu_oflow_irq_0_avs_oflow_writedata -> processor7_0:cpu_oflow_irq_0_avs_oflow_writedata
	wire   [7:0] mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_address;   // mm_interconnect_1:processor7_0_cpu_oflow_irq_0_avs_oflow_address -> processor7_0:cpu_oflow_irq_0_avs_oflow_address
	wire         mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_write;     // mm_interconnect_1:processor7_0_cpu_oflow_irq_0_avs_oflow_write -> processor7_0:cpu_oflow_irq_0_avs_oflow_write
	wire         mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_read;      // mm_interconnect_1:processor7_0_cpu_oflow_irq_0_avs_oflow_read -> processor7_0:cpu_oflow_irq_0_avs_oflow_read
	wire  [31:0] mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_readdata;  // processor7_0:cpu_oflow_irq_0_avs_oflow_readdata -> mm_interconnect_1:processor7_0_cpu_oflow_irq_0_avs_oflow_readdata
	wire  [31:0] mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_writedata; // mm_interconnect_1:processor0_0_cpu_oflow_irq_0_avs_oflow_writedata -> processor0_0:cpu_oflow_irq_0_avs_oflow_writedata
	wire   [7:0] mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_address;   // mm_interconnect_1:processor0_0_cpu_oflow_irq_0_avs_oflow_address -> processor0_0:cpu_oflow_irq_0_avs_oflow_address
	wire         mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_write;     // mm_interconnect_1:processor0_0_cpu_oflow_irq_0_avs_oflow_write -> processor0_0:cpu_oflow_irq_0_avs_oflow_write
	wire         mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_read;      // mm_interconnect_1:processor0_0_cpu_oflow_irq_0_avs_oflow_read -> processor0_0:cpu_oflow_irq_0_avs_oflow_read
	wire  [31:0] mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_readdata;  // processor0_0:cpu_oflow_irq_0_avs_oflow_readdata -> mm_interconnect_1:processor0_0_cpu_oflow_irq_0_avs_oflow_readdata
	wire  [27:0] mm_interconnect_1_processor3_0_dma_0_control_port_slave_writedata;  // mm_interconnect_1:processor3_0_dma_0_control_port_slave_writedata -> processor3_0:dma_0_control_port_slave_writedata
	wire   [2:0] mm_interconnect_1_processor3_0_dma_0_control_port_slave_address;    // mm_interconnect_1:processor3_0_dma_0_control_port_slave_address -> processor3_0:dma_0_control_port_slave_address
	wire         mm_interconnect_1_processor3_0_dma_0_control_port_slave_chipselect; // mm_interconnect_1:processor3_0_dma_0_control_port_slave_chipselect -> processor3_0:dma_0_control_port_slave_chipselect
	wire         mm_interconnect_1_processor3_0_dma_0_control_port_slave_write;      // mm_interconnect_1:processor3_0_dma_0_control_port_slave_write -> processor3_0:dma_0_control_port_slave_write_n
	wire  [27:0] mm_interconnect_1_processor3_0_dma_0_control_port_slave_readdata;   // processor3_0:dma_0_control_port_slave_readdata -> mm_interconnect_1:processor3_0_dma_0_control_port_slave_readdata
	wire  [31:0] mm_interconnect_1_processor7_0_cpu_irq_0_s0_writedata;              // mm_interconnect_1:processor7_0_cpu_irq_0_s0_writedata -> processor7_0:cpu_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processor7_0_cpu_irq_0_s0_address;                // mm_interconnect_1:processor7_0_cpu_irq_0_s0_address -> processor7_0:cpu_irq_0_s0_address
	wire         mm_interconnect_1_processor7_0_cpu_irq_0_s0_write;                  // mm_interconnect_1:processor7_0_cpu_irq_0_s0_write -> processor7_0:cpu_irq_0_s0_write
	wire  [31:0] mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_writedata; // mm_interconnect_1:processor5_0_cpu_oflow_irq_0_avs_oflow_writedata -> processor5_0:cpu_oflow_irq_0_avs_oflow_writedata
	wire   [7:0] mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_address;   // mm_interconnect_1:processor5_0_cpu_oflow_irq_0_avs_oflow_address -> processor5_0:cpu_oflow_irq_0_avs_oflow_address
	wire         mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_write;     // mm_interconnect_1:processor5_0_cpu_oflow_irq_0_avs_oflow_write -> processor5_0:cpu_oflow_irq_0_avs_oflow_write
	wire         mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_read;      // mm_interconnect_1:processor5_0_cpu_oflow_irq_0_avs_oflow_read -> processor5_0:cpu_oflow_irq_0_avs_oflow_read
	wire  [31:0] mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_readdata;  // processor5_0:cpu_oflow_irq_0_avs_oflow_readdata -> mm_interconnect_1:processor5_0_cpu_oflow_irq_0_avs_oflow_readdata
	wire  [31:0] mm_interconnect_1_processor3_0_cpu_irq_0_s0_writedata;              // mm_interconnect_1:processor3_0_cpu_irq_0_s0_writedata -> processor3_0:cpu_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processor3_0_cpu_irq_0_s0_address;                // mm_interconnect_1:processor3_0_cpu_irq_0_s0_address -> processor3_0:cpu_irq_0_s0_address
	wire         mm_interconnect_1_processor3_0_cpu_irq_0_s0_write;                  // mm_interconnect_1:processor3_0_cpu_irq_0_s0_write -> processor3_0:cpu_irq_0_s0_write
	wire  [31:0] mm_interconnect_1_shared_memory_s1_writedata;                       // mm_interconnect_1:shared_memory_s1_writedata -> shared_memory:writedata
	wire   [7:0] mm_interconnect_1_shared_memory_s1_address;                         // mm_interconnect_1:shared_memory_s1_address -> shared_memory:address
	wire         mm_interconnect_1_shared_memory_s1_chipselect;                      // mm_interconnect_1:shared_memory_s1_chipselect -> shared_memory:chipselect
	wire         mm_interconnect_1_shared_memory_s1_clken;                           // mm_interconnect_1:shared_memory_s1_clken -> shared_memory:clken
	wire         mm_interconnect_1_shared_memory_s1_write;                           // mm_interconnect_1:shared_memory_s1_write -> shared_memory:write
	wire  [31:0] mm_interconnect_1_shared_memory_s1_readdata;                        // shared_memory:readdata -> mm_interconnect_1:shared_memory_s1_readdata
	wire   [3:0] mm_interconnect_1_shared_memory_s1_byteenable;                      // mm_interconnect_1:shared_memory_s1_byteenable -> shared_memory:byteenable
	wire  [31:0] mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_writedata; // mm_interconnect_1:processor1_0_cpu_oflow_irq_0_avs_oflow_writedata -> processor1_0:cpu_oflow_irq_0_avs_oflow_writedata
	wire   [7:0] mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_address;   // mm_interconnect_1:processor1_0_cpu_oflow_irq_0_avs_oflow_address -> processor1_0:cpu_oflow_irq_0_avs_oflow_address
	wire         mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_write;     // mm_interconnect_1:processor1_0_cpu_oflow_irq_0_avs_oflow_write -> processor1_0:cpu_oflow_irq_0_avs_oflow_write
	wire         mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_read;      // mm_interconnect_1:processor1_0_cpu_oflow_irq_0_avs_oflow_read -> processor1_0:cpu_oflow_irq_0_avs_oflow_read
	wire  [31:0] mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_readdata;  // processor1_0:cpu_oflow_irq_0_avs_oflow_readdata -> mm_interconnect_1:processor1_0_cpu_oflow_irq_0_avs_oflow_readdata
	wire   [0:0] processor1_0_outgoing_master_burstcount;                            // processor1_0:outgoing_master_burstcount -> mm_interconnect_1:processor1_0_outgoing_master_burstcount
	wire         processor1_0_outgoing_master_waitrequest;                           // mm_interconnect_1:processor1_0_outgoing_master_waitrequest -> processor1_0:outgoing_master_waitrequest
	wire  [26:0] processor1_0_outgoing_master_address;                               // processor1_0:outgoing_master_address -> mm_interconnect_1:processor1_0_outgoing_master_address
	wire  [31:0] processor1_0_outgoing_master_writedata;                             // processor1_0:outgoing_master_writedata -> mm_interconnect_1:processor1_0_outgoing_master_writedata
	wire         processor1_0_outgoing_master_write;                                 // processor1_0:outgoing_master_write -> mm_interconnect_1:processor1_0_outgoing_master_write
	wire         processor1_0_outgoing_master_read;                                  // processor1_0:outgoing_master_read -> mm_interconnect_1:processor1_0_outgoing_master_read
	wire  [31:0] processor1_0_outgoing_master_readdata;                              // mm_interconnect_1:processor1_0_outgoing_master_readdata -> processor1_0:outgoing_master_readdata
	wire         processor1_0_outgoing_master_debugaccess;                           // processor1_0:outgoing_master_debugaccess -> mm_interconnect_1:processor1_0_outgoing_master_debugaccess
	wire   [3:0] processor1_0_outgoing_master_byteenable;                            // processor1_0:outgoing_master_byteenable -> mm_interconnect_1:processor1_0_outgoing_master_byteenable
	wire         processor1_0_outgoing_master_readdatavalid;                         // mm_interconnect_1:processor1_0_outgoing_master_readdatavalid -> processor1_0:outgoing_master_readdatavalid
	wire   [0:0] processorm_0_outgoing_master_burstcount;                            // processorM_0:outgoing_master_burstcount -> mm_interconnect_1:processorM_0_outgoing_master_burstcount
	wire         processorm_0_outgoing_master_waitrequest;                           // mm_interconnect_1:processorM_0_outgoing_master_waitrequest -> processorM_0:outgoing_master_waitrequest
	wire  [26:0] processorm_0_outgoing_master_address;                               // processorM_0:outgoing_master_address -> mm_interconnect_1:processorM_0_outgoing_master_address
	wire  [31:0] processorm_0_outgoing_master_writedata;                             // processorM_0:outgoing_master_writedata -> mm_interconnect_1:processorM_0_outgoing_master_writedata
	wire         processorm_0_outgoing_master_write;                                 // processorM_0:outgoing_master_write -> mm_interconnect_1:processorM_0_outgoing_master_write
	wire         processorm_0_outgoing_master_read;                                  // processorM_0:outgoing_master_read -> mm_interconnect_1:processorM_0_outgoing_master_read
	wire  [31:0] processorm_0_outgoing_master_readdata;                              // mm_interconnect_1:processorM_0_outgoing_master_readdata -> processorM_0:outgoing_master_readdata
	wire         processorm_0_outgoing_master_debugaccess;                           // processorM_0:outgoing_master_debugaccess -> mm_interconnect_1:processorM_0_outgoing_master_debugaccess
	wire   [3:0] processorm_0_outgoing_master_byteenable;                            // processorM_0:outgoing_master_byteenable -> mm_interconnect_1:processorM_0_outgoing_master_byteenable
	wire         processorm_0_outgoing_master_readdatavalid;                         // mm_interconnect_1:processorM_0_outgoing_master_readdatavalid -> processorM_0:outgoing_master_readdatavalid
	wire  [31:0] mm_interconnect_1_processor6_0_cpu_irq_0_s0_writedata;              // mm_interconnect_1:processor6_0_cpu_irq_0_s0_writedata -> processor6_0:cpu_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processor6_0_cpu_irq_0_s0_address;                // mm_interconnect_1:processor6_0_cpu_irq_0_s0_address -> processor6_0:cpu_irq_0_s0_address
	wire         mm_interconnect_1_processor6_0_cpu_irq_0_s0_write;                  // mm_interconnect_1:processor6_0_cpu_irq_0_s0_write -> processor6_0:cpu_irq_0_s0_write
	wire         processor6_0_fingerprint_0_avalon_master_waitrequest;               // mm_interconnect_1:processor6_0_fingerprint_0_avalon_master_waitrequest -> processor6_0:fingerprint_0_avalon_master_waitrequest
	wire  [26:0] processor6_0_fingerprint_0_avalon_master_address;                   // processor6_0:fingerprint_0_avalon_master_address -> mm_interconnect_1:processor6_0_fingerprint_0_avalon_master_address
	wire  [31:0] processor6_0_fingerprint_0_avalon_master_writedata;                 // processor6_0:fingerprint_0_avalon_master_writedata -> mm_interconnect_1:processor6_0_fingerprint_0_avalon_master_writedata
	wire         processor6_0_fingerprint_0_avalon_master_write;                     // processor6_0:fingerprint_0_avalon_master_write -> mm_interconnect_1:processor6_0_fingerprint_0_avalon_master_write
	wire         processor6_0_fingerprint_0_avalon_master_read;                      // processor6_0:fingerprint_0_avalon_master_read -> mm_interconnect_1:processor6_0_fingerprint_0_avalon_master_read
	wire  [31:0] processor6_0_fingerprint_0_avalon_master_readdata;                  // mm_interconnect_1:processor6_0_fingerprint_0_avalon_master_readdata -> processor6_0:fingerprint_0_avalon_master_readdata
	wire  [31:0] mm_interconnect_1_mutex_0_s1_writedata;                             // mm_interconnect_1:mutex_0_s1_writedata -> mutex_0:data_from_cpu
	wire   [0:0] mm_interconnect_1_mutex_0_s1_address;                               // mm_interconnect_1:mutex_0_s1_address -> mutex_0:address
	wire         mm_interconnect_1_mutex_0_s1_chipselect;                            // mm_interconnect_1:mutex_0_s1_chipselect -> mutex_0:chipselect
	wire         mm_interconnect_1_mutex_0_s1_write;                                 // mm_interconnect_1:mutex_0_s1_write -> mutex_0:write
	wire         mm_interconnect_1_mutex_0_s1_read;                                  // mm_interconnect_1:mutex_0_s1_read -> mutex_0:read
	wire  [31:0] mm_interconnect_1_mutex_0_s1_readdata;                              // mutex_0:data_to_cpu -> mm_interconnect_1:mutex_0_s1_readdata
	wire  [31:0] mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_writedata; // mm_interconnect_1:processor3_0_cpu_oflow_irq_0_avs_oflow_writedata -> processor3_0:cpu_oflow_irq_0_avs_oflow_writedata
	wire   [7:0] mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_address;   // mm_interconnect_1:processor3_0_cpu_oflow_irq_0_avs_oflow_address -> processor3_0:cpu_oflow_irq_0_avs_oflow_address
	wire         mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_write;     // mm_interconnect_1:processor3_0_cpu_oflow_irq_0_avs_oflow_write -> processor3_0:cpu_oflow_irq_0_avs_oflow_write
	wire         mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_read;      // mm_interconnect_1:processor3_0_cpu_oflow_irq_0_avs_oflow_read -> processor3_0:cpu_oflow_irq_0_avs_oflow_read
	wire  [31:0] mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_readdata;  // processor3_0:cpu_oflow_irq_0_avs_oflow_readdata -> mm_interconnect_1:processor3_0_cpu_oflow_irq_0_avs_oflow_readdata
	wire   [0:0] processor7_0_out_system_bridge_m0_burstcount;                       // processor7_0:out_system_bridge_m0_burstcount -> mm_interconnect_1:processor7_0_out_system_bridge_m0_burstcount
	wire         processor7_0_out_system_bridge_m0_waitrequest;                      // mm_interconnect_1:processor7_0_out_system_bridge_m0_waitrequest -> processor7_0:out_system_bridge_m0_waitrequest
	wire  [26:0] processor7_0_out_system_bridge_m0_address;                          // processor7_0:out_system_bridge_m0_address -> mm_interconnect_1:processor7_0_out_system_bridge_m0_address
	wire  [31:0] processor7_0_out_system_bridge_m0_writedata;                        // processor7_0:out_system_bridge_m0_writedata -> mm_interconnect_1:processor7_0_out_system_bridge_m0_writedata
	wire         processor7_0_out_system_bridge_m0_write;                            // processor7_0:out_system_bridge_m0_write -> mm_interconnect_1:processor7_0_out_system_bridge_m0_write
	wire         processor7_0_out_system_bridge_m0_read;                             // processor7_0:out_system_bridge_m0_read -> mm_interconnect_1:processor7_0_out_system_bridge_m0_read
	wire  [31:0] processor7_0_out_system_bridge_m0_readdata;                         // mm_interconnect_1:processor7_0_out_system_bridge_m0_readdata -> processor7_0:out_system_bridge_m0_readdata
	wire         processor7_0_out_system_bridge_m0_debugaccess;                      // processor7_0:out_system_bridge_m0_debugaccess -> mm_interconnect_1:processor7_0_out_system_bridge_m0_debugaccess
	wire   [3:0] processor7_0_out_system_bridge_m0_byteenable;                       // processor7_0:out_system_bridge_m0_byteenable -> mm_interconnect_1:processor7_0_out_system_bridge_m0_byteenable
	wire         processor7_0_out_system_bridge_m0_readdatavalid;                    // mm_interconnect_1:processor7_0_out_system_bridge_m0_readdatavalid -> processor7_0:out_system_bridge_m0_readdatavalid
	wire  [27:0] mm_interconnect_1_processor1_0_dma_0_control_port_slave_writedata;  // mm_interconnect_1:processor1_0_dma_0_control_port_slave_writedata -> processor1_0:dma_0_control_port_slave_writedata
	wire   [2:0] mm_interconnect_1_processor1_0_dma_0_control_port_slave_address;    // mm_interconnect_1:processor1_0_dma_0_control_port_slave_address -> processor1_0:dma_0_control_port_slave_address
	wire         mm_interconnect_1_processor1_0_dma_0_control_port_slave_chipselect; // mm_interconnect_1:processor1_0_dma_0_control_port_slave_chipselect -> processor1_0:dma_0_control_port_slave_chipselect
	wire         mm_interconnect_1_processor1_0_dma_0_control_port_slave_write;      // mm_interconnect_1:processor1_0_dma_0_control_port_slave_write -> processor1_0:dma_0_control_port_slave_write_n
	wire  [27:0] mm_interconnect_1_processor1_0_dma_0_control_port_slave_readdata;   // processor1_0:dma_0_control_port_slave_readdata -> mm_interconnect_1:processor1_0_dma_0_control_port_slave_readdata
	wire  [27:0] mm_interconnect_1_processor7_0_dma_0_control_port_slave_writedata;  // mm_interconnect_1:processor7_0_dma_0_control_port_slave_writedata -> processor7_0:dma_0_control_port_slave_writedata
	wire   [2:0] mm_interconnect_1_processor7_0_dma_0_control_port_slave_address;    // mm_interconnect_1:processor7_0_dma_0_control_port_slave_address -> processor7_0:dma_0_control_port_slave_address
	wire         mm_interconnect_1_processor7_0_dma_0_control_port_slave_chipselect; // mm_interconnect_1:processor7_0_dma_0_control_port_slave_chipselect -> processor7_0:dma_0_control_port_slave_chipselect
	wire         mm_interconnect_1_processor7_0_dma_0_control_port_slave_write;      // mm_interconnect_1:processor7_0_dma_0_control_port_slave_write -> processor7_0:dma_0_control_port_slave_write_n
	wire  [27:0] mm_interconnect_1_processor7_0_dma_0_control_port_slave_readdata;   // processor7_0:dma_0_control_port_slave_readdata -> mm_interconnect_1:processor7_0_dma_0_control_port_slave_readdata
	wire  [27:0] mm_interconnect_1_processor4_0_dma_0_control_port_slave_writedata;  // mm_interconnect_1:processor4_0_dma_0_control_port_slave_writedata -> processor4_0:dma_0_control_port_slave_writedata
	wire   [2:0] mm_interconnect_1_processor4_0_dma_0_control_port_slave_address;    // mm_interconnect_1:processor4_0_dma_0_control_port_slave_address -> processor4_0:dma_0_control_port_slave_address
	wire         mm_interconnect_1_processor4_0_dma_0_control_port_slave_chipselect; // mm_interconnect_1:processor4_0_dma_0_control_port_slave_chipselect -> processor4_0:dma_0_control_port_slave_chipselect
	wire         mm_interconnect_1_processor4_0_dma_0_control_port_slave_write;      // mm_interconnect_1:processor4_0_dma_0_control_port_slave_write -> processor4_0:dma_0_control_port_slave_write_n
	wire  [27:0] mm_interconnect_1_processor4_0_dma_0_control_port_slave_readdata;   // processor4_0:dma_0_control_port_slave_readdata -> mm_interconnect_1:processor4_0_dma_0_control_port_slave_readdata
	wire   [0:0] processor3_0_out_system_bridge_m0_burstcount;                       // processor3_0:out_system_bridge_m0_burstcount -> mm_interconnect_1:processor3_0_out_system_bridge_m0_burstcount
	wire         processor3_0_out_system_bridge_m0_waitrequest;                      // mm_interconnect_1:processor3_0_out_system_bridge_m0_waitrequest -> processor3_0:out_system_bridge_m0_waitrequest
	wire  [26:0] processor3_0_out_system_bridge_m0_address;                          // processor3_0:out_system_bridge_m0_address -> mm_interconnect_1:processor3_0_out_system_bridge_m0_address
	wire  [31:0] processor3_0_out_system_bridge_m0_writedata;                        // processor3_0:out_system_bridge_m0_writedata -> mm_interconnect_1:processor3_0_out_system_bridge_m0_writedata
	wire         processor3_0_out_system_bridge_m0_write;                            // processor3_0:out_system_bridge_m0_write -> mm_interconnect_1:processor3_0_out_system_bridge_m0_write
	wire         processor3_0_out_system_bridge_m0_read;                             // processor3_0:out_system_bridge_m0_read -> mm_interconnect_1:processor3_0_out_system_bridge_m0_read
	wire  [31:0] processor3_0_out_system_bridge_m0_readdata;                         // mm_interconnect_1:processor3_0_out_system_bridge_m0_readdata -> processor3_0:out_system_bridge_m0_readdata
	wire         processor3_0_out_system_bridge_m0_debugaccess;                      // processor3_0:out_system_bridge_m0_debugaccess -> mm_interconnect_1:processor3_0_out_system_bridge_m0_debugaccess
	wire   [3:0] processor3_0_out_system_bridge_m0_byteenable;                       // processor3_0:out_system_bridge_m0_byteenable -> mm_interconnect_1:processor3_0_out_system_bridge_m0_byteenable
	wire         processor3_0_out_system_bridge_m0_readdatavalid;                    // mm_interconnect_1:processor3_0_out_system_bridge_m0_readdatavalid -> processor3_0:out_system_bridge_m0_readdatavalid
	wire  [31:0] mm_interconnect_1_processorm_0_cpu_irq_0_s0_writedata;              // mm_interconnect_1:processorM_0_cpu_irq_0_s0_writedata -> processorM_0:cpu_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processorm_0_cpu_irq_0_s0_address;                // mm_interconnect_1:processorM_0_cpu_irq_0_s0_address -> processorM_0:cpu_irq_0_s0_address
	wire         mm_interconnect_1_processorm_0_cpu_irq_0_s0_write;                  // mm_interconnect_1:processorM_0_cpu_irq_0_s0_write -> processorM_0:cpu_irq_0_s0_write
	wire         cfpu_0_oflow_waitrequest;                                           // mm_interconnect_1:cfpu_0_oflow_waitrequest -> cfpu_0:oflow_waitrequest
	wire  [26:0] cfpu_0_oflow_address;                                               // cfpu_0:oflow_address -> mm_interconnect_1:cfpu_0_oflow_address
	wire  [31:0] cfpu_0_oflow_writedata;                                             // cfpu_0:oflow_writedata -> mm_interconnect_1:cfpu_0_oflow_writedata
	wire         cfpu_0_oflow_write;                                                 // cfpu_0:oflow_write -> mm_interconnect_1:cfpu_0_oflow_write
	wire         processor5_0_fingerprint_0_avalon_master_waitrequest;               // mm_interconnect_1:processor5_0_fingerprint_0_avalon_master_waitrequest -> processor5_0:fingerprint_0_avalon_master_waitrequest
	wire  [26:0] processor5_0_fingerprint_0_avalon_master_address;                   // processor5_0:fingerprint_0_avalon_master_address -> mm_interconnect_1:processor5_0_fingerprint_0_avalon_master_address
	wire  [31:0] processor5_0_fingerprint_0_avalon_master_writedata;                 // processor5_0:fingerprint_0_avalon_master_writedata -> mm_interconnect_1:processor5_0_fingerprint_0_avalon_master_writedata
	wire         processor5_0_fingerprint_0_avalon_master_write;                     // processor5_0:fingerprint_0_avalon_master_write -> mm_interconnect_1:processor5_0_fingerprint_0_avalon_master_write
	wire         processor5_0_fingerprint_0_avalon_master_read;                      // processor5_0:fingerprint_0_avalon_master_read -> mm_interconnect_1:processor5_0_fingerprint_0_avalon_master_read
	wire  [31:0] processor5_0_fingerprint_0_avalon_master_readdata;                  // mm_interconnect_1:processor5_0_fingerprint_0_avalon_master_readdata -> processor5_0:fingerprint_0_avalon_master_readdata
	wire  [27:0] mm_interconnect_1_processor0_0_dma_0_control_port_slave_writedata;  // mm_interconnect_1:processor0_0_dma_0_control_port_slave_writedata -> processor0_0:dma_0_control_port_slave_writedata
	wire   [2:0] mm_interconnect_1_processor0_0_dma_0_control_port_slave_address;    // mm_interconnect_1:processor0_0_dma_0_control_port_slave_address -> processor0_0:dma_0_control_port_slave_address
	wire         mm_interconnect_1_processor0_0_dma_0_control_port_slave_chipselect; // mm_interconnect_1:processor0_0_dma_0_control_port_slave_chipselect -> processor0_0:dma_0_control_port_slave_chipselect
	wire         mm_interconnect_1_processor0_0_dma_0_control_port_slave_write;      // mm_interconnect_1:processor0_0_dma_0_control_port_slave_write -> processor0_0:dma_0_control_port_slave_write_n
	wire  [27:0] mm_interconnect_1_processor0_0_dma_0_control_port_slave_readdata;   // processor0_0:dma_0_control_port_slave_readdata -> mm_interconnect_1:processor0_0_dma_0_control_port_slave_readdata
	wire   [0:0] processor5_0_out_system_bridge_m0_burstcount;                       // processor5_0:out_system_bridge_m0_burstcount -> mm_interconnect_1:processor5_0_out_system_bridge_m0_burstcount
	wire         processor5_0_out_system_bridge_m0_waitrequest;                      // mm_interconnect_1:processor5_0_out_system_bridge_m0_waitrequest -> processor5_0:out_system_bridge_m0_waitrequest
	wire  [26:0] processor5_0_out_system_bridge_m0_address;                          // processor5_0:out_system_bridge_m0_address -> mm_interconnect_1:processor5_0_out_system_bridge_m0_address
	wire  [31:0] processor5_0_out_system_bridge_m0_writedata;                        // processor5_0:out_system_bridge_m0_writedata -> mm_interconnect_1:processor5_0_out_system_bridge_m0_writedata
	wire         processor5_0_out_system_bridge_m0_write;                            // processor5_0:out_system_bridge_m0_write -> mm_interconnect_1:processor5_0_out_system_bridge_m0_write
	wire         processor5_0_out_system_bridge_m0_read;                             // processor5_0:out_system_bridge_m0_read -> mm_interconnect_1:processor5_0_out_system_bridge_m0_read
	wire  [31:0] processor5_0_out_system_bridge_m0_readdata;                         // mm_interconnect_1:processor5_0_out_system_bridge_m0_readdata -> processor5_0:out_system_bridge_m0_readdata
	wire         processor5_0_out_system_bridge_m0_debugaccess;                      // processor5_0:out_system_bridge_m0_debugaccess -> mm_interconnect_1:processor5_0_out_system_bridge_m0_debugaccess
	wire   [3:0] processor5_0_out_system_bridge_m0_byteenable;                       // processor5_0:out_system_bridge_m0_byteenable -> mm_interconnect_1:processor5_0_out_system_bridge_m0_byteenable
	wire         processor5_0_out_system_bridge_m0_readdatavalid;                    // mm_interconnect_1:processor5_0_out_system_bridge_m0_readdatavalid -> processor5_0:out_system_bridge_m0_readdatavalid
	wire         processor0_0_fingerprint_0_avalon_master_waitrequest;               // mm_interconnect_1:processor0_0_fingerprint_0_avalon_master_waitrequest -> processor0_0:fingerprint_0_avalon_master_waitrequest
	wire  [26:0] processor0_0_fingerprint_0_avalon_master_address;                   // processor0_0:fingerprint_0_avalon_master_address -> mm_interconnect_1:processor0_0_fingerprint_0_avalon_master_address
	wire  [31:0] processor0_0_fingerprint_0_avalon_master_writedata;                 // processor0_0:fingerprint_0_avalon_master_writedata -> mm_interconnect_1:processor0_0_fingerprint_0_avalon_master_writedata
	wire         processor0_0_fingerprint_0_avalon_master_write;                     // processor0_0:fingerprint_0_avalon_master_write -> mm_interconnect_1:processor0_0_fingerprint_0_avalon_master_write
	wire         processor0_0_fingerprint_0_avalon_master_read;                      // processor0_0:fingerprint_0_avalon_master_read -> mm_interconnect_1:processor0_0_fingerprint_0_avalon_master_read
	wire  [31:0] processor0_0_fingerprint_0_avalon_master_readdata;                  // mm_interconnect_1:processor0_0_fingerprint_0_avalon_master_readdata -> processor0_0:fingerprint_0_avalon_master_readdata
	wire  [31:0] mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_writedata; // mm_interconnect_1:processor4_0_cpu_oflow_irq_0_avs_oflow_writedata -> processor4_0:cpu_oflow_irq_0_avs_oflow_writedata
	wire   [7:0] mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_address;   // mm_interconnect_1:processor4_0_cpu_oflow_irq_0_avs_oflow_address -> processor4_0:cpu_oflow_irq_0_avs_oflow_address
	wire         mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_write;     // mm_interconnect_1:processor4_0_cpu_oflow_irq_0_avs_oflow_write -> processor4_0:cpu_oflow_irq_0_avs_oflow_write
	wire         mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_read;      // mm_interconnect_1:processor4_0_cpu_oflow_irq_0_avs_oflow_read -> processor4_0:cpu_oflow_irq_0_avs_oflow_read
	wire  [31:0] mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_readdata;  // processor4_0:cpu_oflow_irq_0_avs_oflow_readdata -> mm_interconnect_1:processor4_0_cpu_oflow_irq_0_avs_oflow_readdata
	wire         processor1_0_fingerprint_0_avalon_master_waitrequest;               // mm_interconnect_1:processor1_0_fingerprint_0_avalon_master_waitrequest -> processor1_0:fingerprint_0_avalon_master_waitrequest
	wire  [26:0] processor1_0_fingerprint_0_avalon_master_address;                   // processor1_0:fingerprint_0_avalon_master_address -> mm_interconnect_1:processor1_0_fingerprint_0_avalon_master_address
	wire  [31:0] processor1_0_fingerprint_0_avalon_master_writedata;                 // processor1_0:fingerprint_0_avalon_master_writedata -> mm_interconnect_1:processor1_0_fingerprint_0_avalon_master_writedata
	wire         processor1_0_fingerprint_0_avalon_master_write;                     // processor1_0:fingerprint_0_avalon_master_write -> mm_interconnect_1:processor1_0_fingerprint_0_avalon_master_write
	wire         processor1_0_fingerprint_0_avalon_master_read;                      // processor1_0:fingerprint_0_avalon_master_read -> mm_interconnect_1:processor1_0_fingerprint_0_avalon_master_read
	wire  [31:0] processor1_0_fingerprint_0_avalon_master_readdata;                  // mm_interconnect_1:processor1_0_fingerprint_0_avalon_master_readdata -> processor1_0:fingerprint_0_avalon_master_readdata
	wire         processor7_0_fingerprint_0_avalon_master_waitrequest;               // mm_interconnect_1:processor7_0_fingerprint_0_avalon_master_waitrequest -> processor7_0:fingerprint_0_avalon_master_waitrequest
	wire  [26:0] processor7_0_fingerprint_0_avalon_master_address;                   // processor7_0:fingerprint_0_avalon_master_address -> mm_interconnect_1:processor7_0_fingerprint_0_avalon_master_address
	wire  [31:0] processor7_0_fingerprint_0_avalon_master_writedata;                 // processor7_0:fingerprint_0_avalon_master_writedata -> mm_interconnect_1:processor7_0_fingerprint_0_avalon_master_writedata
	wire         processor7_0_fingerprint_0_avalon_master_write;                     // processor7_0:fingerprint_0_avalon_master_write -> mm_interconnect_1:processor7_0_fingerprint_0_avalon_master_write
	wire         processor7_0_fingerprint_0_avalon_master_read;                      // processor7_0:fingerprint_0_avalon_master_read -> mm_interconnect_1:processor7_0_fingerprint_0_avalon_master_read
	wire  [31:0] processor7_0_fingerprint_0_avalon_master_readdata;                  // mm_interconnect_1:processor7_0_fingerprint_0_avalon_master_readdata -> processor7_0:fingerprint_0_avalon_master_readdata
	wire  [31:0] mm_interconnect_1_memory_0_memory_delay_0_csr_writedata;            // mm_interconnect_1:memory_0_memory_delay_0_csr_writedata -> memory_0:memory_delay_0_csr_writedata
	wire   [2:0] mm_interconnect_1_memory_0_memory_delay_0_csr_address;              // mm_interconnect_1:memory_0_memory_delay_0_csr_address -> memory_0:memory_delay_0_csr_address
	wire         mm_interconnect_1_memory_0_memory_delay_0_csr_write;                // mm_interconnect_1:memory_0_memory_delay_0_csr_write -> memory_0:memory_delay_0_csr_write
	wire  [31:0] mm_interconnect_1_processor0_0_cpu_irq_0_s0_writedata;              // mm_interconnect_1:processor0_0_cpu_irq_0_s0_writedata -> processor0_0:cpu_irq_0_s0_writedata
	wire   [7:0] mm_interconnect_1_processor0_0_cpu_irq_0_s0_address;                // mm_interconnect_1:processor0_0_cpu_irq_0_s0_address -> processor0_0:cpu_irq_0_s0_address
	wire         mm_interconnect_1_processor0_0_cpu_irq_0_s0_write;                  // mm_interconnect_1:processor0_0_cpu_irq_0_s0_write -> processor0_0:cpu_irq_0_s0_write
	wire   [0:0] processor4_0_out_system_bridge_m0_burstcount;                       // processor4_0:out_system_bridge_m0_burstcount -> mm_interconnect_1:processor4_0_out_system_bridge_m0_burstcount
	wire         processor4_0_out_system_bridge_m0_waitrequest;                      // mm_interconnect_1:processor4_0_out_system_bridge_m0_waitrequest -> processor4_0:out_system_bridge_m0_waitrequest
	wire  [26:0] processor4_0_out_system_bridge_m0_address;                          // processor4_0:out_system_bridge_m0_address -> mm_interconnect_1:processor4_0_out_system_bridge_m0_address
	wire  [31:0] processor4_0_out_system_bridge_m0_writedata;                        // processor4_0:out_system_bridge_m0_writedata -> mm_interconnect_1:processor4_0_out_system_bridge_m0_writedata
	wire         processor4_0_out_system_bridge_m0_write;                            // processor4_0:out_system_bridge_m0_write -> mm_interconnect_1:processor4_0_out_system_bridge_m0_write
	wire         processor4_0_out_system_bridge_m0_read;                             // processor4_0:out_system_bridge_m0_read -> mm_interconnect_1:processor4_0_out_system_bridge_m0_read
	wire  [31:0] processor4_0_out_system_bridge_m0_readdata;                         // mm_interconnect_1:processor4_0_out_system_bridge_m0_readdata -> processor4_0:out_system_bridge_m0_readdata
	wire         processor4_0_out_system_bridge_m0_debugaccess;                      // processor4_0:out_system_bridge_m0_debugaccess -> mm_interconnect_1:processor4_0_out_system_bridge_m0_debugaccess
	wire   [3:0] processor4_0_out_system_bridge_m0_byteenable;                       // processor4_0:out_system_bridge_m0_byteenable -> mm_interconnect_1:processor4_0_out_system_bridge_m0_byteenable
	wire         processor4_0_out_system_bridge_m0_readdatavalid;                    // mm_interconnect_1:processor4_0_out_system_bridge_m0_readdatavalid -> processor4_0:out_system_bridge_m0_readdatavalid
	wire         processor4_0_fingerprint_0_avalon_master_waitrequest;               // mm_interconnect_1:processor4_0_fingerprint_0_avalon_master_waitrequest -> processor4_0:fingerprint_0_avalon_master_waitrequest
	wire  [26:0] processor4_0_fingerprint_0_avalon_master_address;                   // processor4_0:fingerprint_0_avalon_master_address -> mm_interconnect_1:processor4_0_fingerprint_0_avalon_master_address
	wire  [31:0] processor4_0_fingerprint_0_avalon_master_writedata;                 // processor4_0:fingerprint_0_avalon_master_writedata -> mm_interconnect_1:processor4_0_fingerprint_0_avalon_master_writedata
	wire         processor4_0_fingerprint_0_avalon_master_write;                     // processor4_0:fingerprint_0_avalon_master_write -> mm_interconnect_1:processor4_0_fingerprint_0_avalon_master_write
	wire         processor4_0_fingerprint_0_avalon_master_read;                      // processor4_0:fingerprint_0_avalon_master_read -> mm_interconnect_1:processor4_0_fingerprint_0_avalon_master_read
	wire  [31:0] processor4_0_fingerprint_0_avalon_master_readdata;                  // mm_interconnect_1:processor4_0_fingerprint_0_avalon_master_readdata -> processor4_0:fingerprint_0_avalon_master_readdata
	wire         irq_mapper_receiver0_irq;                                           // processor0_0:dma_0_irq_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                           // processor1_0:dma_0_irq_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                           // processor2_0:dma_0_irq_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                           // processor3_0:dma_0_irq_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                           // processor4_0:dma_0_irq_irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                           // processor5_0:dma_0_irq_irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                           // processor6_0:dma_0_irq_irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                           // processor7_0:dma_0_irq_irq -> irq_mapper:receiver7_irq
	wire   [7:0] processorm_0_dma_0_irq_receiver_irq_irq;                            // irq_mapper:sender_irq -> processorM_0:dma_0_irq_receiver_irq_irq
	wire         rst_controller_reset_out_reset;                                     // rst_controller:reset_out -> [cfpu_0:reset, irq_mapper:reset, mm_bridge_0:reset, mm_interconnect_0:memory_0_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mm_bridge_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:cfpu_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:processor1_0_reset_reset_bridge_in_reset_reset, mutex_0:reset_n, rst_translator:in_reset, shared_memory:reset, sys_id:reset_n]
	wire         rst_controller_reset_out_reset_req;                                 // rst_controller:reset_req -> [rst_translator:reset_req_in, shared_memory:reset_req]

	nios_fprint_sys_id sys_id (
		.clock    (clk_clk),                                         //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	nios_fprint_shared_memory shared_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_1_shared_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_1_shared_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_1_shared_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_1_shared_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_1_shared_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_1_shared_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_1_shared_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)             //       .reset_req
	);

	nios_fprint_mutex_0 mutex_0 (
		.reset_n       (~rst_controller_reset_out_reset),         // reset.reset_n
		.clk           (clk_clk),                                 //   clk.clk
		.chipselect    (mm_interconnect_1_mutex_0_s1_chipselect), //    s1.chipselect
		.data_from_cpu (mm_interconnect_1_mutex_0_s1_writedata),  //      .writedata
		.read          (mm_interconnect_1_mutex_0_s1_read),       //      .read
		.write         (mm_interconnect_1_mutex_0_s1_write),      //      .write
		.data_to_cpu   (mm_interconnect_1_mutex_0_s1_readdata),   //      .readdata
		.address       (mm_interconnect_1_mutex_0_s1_address)     //      .address
	);

	cfpu cfpu_0 (
		.clk                (clk_clk),                                     //  clock.clk
		.reset              (rst_controller_reset_out_reset),              //  reset.reset
		.csr_address        (mm_interconnect_1_cfpu_0_csr_address),        //    csr.address
		.csr_read           (mm_interconnect_1_cfpu_0_csr_read),           //       .read
		.csr_readdata       (mm_interconnect_1_cfpu_0_csr_readdata),       //       .readdata
		.csr_write          (mm_interconnect_1_cfpu_0_csr_write),          //       .write
		.csr_writedata      (mm_interconnect_1_cfpu_0_csr_writedata),      //       .writedata
		.csr_waitrequest    (mm_interconnect_1_cfpu_0_csr_waitrequest),    //       .waitrequest
		.fprint_address     (mm_interconnect_0_cfpu_0_fprint_address),     // fprint.address
		.fprint_write       (mm_interconnect_0_cfpu_0_fprint_write),       //       .write
		.fprint_writedata   (mm_interconnect_0_cfpu_0_fprint_writedata),   //       .writedata
		.fprint_waitrequest (mm_interconnect_0_cfpu_0_fprint_waitrequest), //       .waitrequest
		.oflow_write        (cfpu_0_oflow_write),                          //  oflow.write
		.oflow_writedata    (cfpu_0_oflow_writedata),                      //       .writedata
		.oflow_address      (cfpu_0_oflow_address),                        //       .address
		.oflow_waitrequest  (cfpu_0_oflow_waitrequest),                    //       .waitrequest
		.irq                (cfpu_0_irq_export)                            //    irq.export
	);

	nios_fprint_memory_0 memory_0 (
		.clk_clk                      (clk_clk),                                                 //                clk.clk
		.reset_reset_n                (reset_reset_n),                                           //              reset.reset_n
		.mm_bridge_0_s0_waitrequest   (mm_interconnect_0_memory_0_mm_bridge_0_s0_waitrequest),   //     mm_bridge_0_s0.waitrequest
		.mm_bridge_0_s0_readdata      (mm_interconnect_0_memory_0_mm_bridge_0_s0_readdata),      //                   .readdata
		.mm_bridge_0_s0_readdatavalid (mm_interconnect_0_memory_0_mm_bridge_0_s0_readdatavalid), //                   .readdatavalid
		.mm_bridge_0_s0_burstcount    (mm_interconnect_0_memory_0_mm_bridge_0_s0_burstcount),    //                   .burstcount
		.mm_bridge_0_s0_writedata     (mm_interconnect_0_memory_0_mm_bridge_0_s0_writedata),     //                   .writedata
		.mm_bridge_0_s0_address       (mm_interconnect_0_memory_0_mm_bridge_0_s0_address),       //                   .address
		.mm_bridge_0_s0_write         (mm_interconnect_0_memory_0_mm_bridge_0_s0_write),         //                   .write
		.mm_bridge_0_s0_read          (mm_interconnect_0_memory_0_mm_bridge_0_s0_read),          //                   .read
		.mm_bridge_0_s0_byteenable    (mm_interconnect_0_memory_0_mm_bridge_0_s0_byteenable),    //                   .byteenable
		.mm_bridge_0_s0_debugaccess   (mm_interconnect_0_memory_0_mm_bridge_0_s0_debugaccess),   //                   .debugaccess
		.memory_delay_0_csr_address   (mm_interconnect_1_memory_0_memory_delay_0_csr_address),   // memory_delay_0_csr.address
		.memory_delay_0_csr_write     (mm_interconnect_1_memory_0_memory_delay_0_csr_write),     //                   .write
		.memory_delay_0_csr_writedata (mm_interconnect_1_memory_0_memory_delay_0_csr_writedata)  //                   .writedata
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (25),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge_0 (
		.clk              (clk_clk),                                        //   clk.clk
		.reset            (rst_controller_reset_out_reset),                 // reset.reset
		.s0_waitrequest   (mm_interconnect_1_mm_bridge_0_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_1_mm_bridge_0_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_1_mm_bridge_0_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_1_mm_bridge_0_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_1_mm_bridge_0_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_1_mm_bridge_0_s0_address),       //      .address
		.s0_write         (mm_interconnect_1_mm_bridge_0_s0_write),         //      .write
		.s0_read          (mm_interconnect_1_mm_bridge_0_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_1_mm_bridge_0_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_1_mm_bridge_0_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (mm_bridge_0_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (mm_bridge_0_m0_readdata),                        //      .readdata
		.m0_readdatavalid (mm_bridge_0_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (mm_bridge_0_m0_burstcount),                      //      .burstcount
		.m0_writedata     (mm_bridge_0_m0_writedata),                       //      .writedata
		.m0_address       (mm_bridge_0_m0_address),                         //      .address
		.m0_write         (mm_bridge_0_m0_write),                           //      .write
		.m0_read          (mm_bridge_0_m0_read),                            //      .read
		.m0_byteenable    (mm_bridge_0_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (mm_bridge_0_m0_debugaccess)                      //      .debugaccess
	);

	nios_fprint_processor1_0 processor1_0 (
		.philosopher_clk_in_clk                  (clk_clk),                                                            //             philosopher_clk_in.clk
		.outgoing_master_waitrequest             (processor1_0_outgoing_master_waitrequest),                           //                outgoing_master.waitrequest
		.outgoing_master_readdata                (processor1_0_outgoing_master_readdata),                              //                               .readdata
		.outgoing_master_readdatavalid           (processor1_0_outgoing_master_readdatavalid),                         //                               .readdatavalid
		.outgoing_master_burstcount              (processor1_0_outgoing_master_burstcount),                            //                               .burstcount
		.outgoing_master_writedata               (processor1_0_outgoing_master_writedata),                             //                               .writedata
		.outgoing_master_address                 (processor1_0_outgoing_master_address),                               //                               .address
		.outgoing_master_write                   (processor1_0_outgoing_master_write),                                 //                               .write
		.outgoing_master_read                    (processor1_0_outgoing_master_read),                                  //                               .read
		.outgoing_master_byteenable              (processor1_0_outgoing_master_byteenable),                            //                               .byteenable
		.outgoing_master_debugaccess             (processor1_0_outgoing_master_debugaccess),                           //                               .debugaccess
		.button_pio_external_connection_export   (),                                                                   // button_pio_external_connection.export
		.reset_reset_n                           (reset_reset_n),                                                      //                          reset.reset_n
		.cpu1_jtag_debug_module_reset_reset      (),                                                                   //   cpu1_jtag_debug_module_reset.reset
		.cpu1_irq_0_s0_address                   (mm_interconnect_1_processor1_0_cpu1_irq_0_s0_address),               //                  cpu1_irq_0_s0.address
		.cpu1_irq_0_s0_write                     (mm_interconnect_1_processor1_0_cpu1_irq_0_s0_write),                 //                               .write
		.cpu1_irq_0_s0_writedata                 (mm_interconnect_1_processor1_0_cpu1_irq_0_s0_writedata),             //                               .writedata
		.dma_0_control_port_slave_address        (mm_interconnect_1_processor1_0_dma_0_control_port_slave_address),    //       dma_0_control_port_slave.address
		.dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor1_0_dma_0_control_port_slave_chipselect), //                               .chipselect
		.dma_0_control_port_slave_readdata       (mm_interconnect_1_processor1_0_dma_0_control_port_slave_readdata),   //                               .readdata
		.dma_0_control_port_slave_write_n        (~mm_interconnect_1_processor1_0_dma_0_control_port_slave_write),     //                               .write_n
		.dma_0_control_port_slave_writedata      (mm_interconnect_1_processor1_0_dma_0_control_port_slave_writedata),  //                               .writedata
		.dma_0_irq_irq                           (irq_mapper_receiver1_irq),                                           //                      dma_0_irq.irq
		.fingerprint_0_avalon_master_writedata   (processor1_0_fingerprint_0_avalon_master_writedata),                 //    fingerprint_0_avalon_master.writedata
		.fingerprint_0_avalon_master_write       (processor1_0_fingerprint_0_avalon_master_write),                     //                               .write
		.fingerprint_0_avalon_master_readdata    (processor1_0_fingerprint_0_avalon_master_readdata),                  //                               .readdata
		.fingerprint_0_avalon_master_waitrequest (processor1_0_fingerprint_0_avalon_master_waitrequest),               //                               .waitrequest
		.fingerprint_0_avalon_master_read        (processor1_0_fingerprint_0_avalon_master_read),                      //                               .read
		.fingerprint_0_avalon_master_address     (processor1_0_fingerprint_0_avalon_master_address),                   //                               .address
		.cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_address),   //      cpu_oflow_irq_0_avs_oflow.address
		.cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_write),     //                               .write
		.cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_writedata), //                               .writedata
		.cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_read),      //                               .read
		.cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_readdata)   //                               .readdata
	);

	nios_fprint_processor0_0 processor0_0 (
		.philosopher_clk_in_clk                  (clk_clk),                                                            //             philosopher_clk_in.clk
		.button_pio_external_connection_export   (),                                                                   // button_pio_external_connection.export
		.cpu0_jtag_debug_module_reset_reset      (),                                                                   //   cpu0_jtag_debug_module_reset.reset
		.reset_reset_n                           (reset_reset_n),                                                      //                          reset.reset_n
		.cpu_irq_0_s0_address                    (mm_interconnect_1_processor0_0_cpu_irq_0_s0_address),                //                   cpu_irq_0_s0.address
		.cpu_irq_0_s0_write                      (mm_interconnect_1_processor0_0_cpu_irq_0_s0_write),                  //                               .write
		.cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor0_0_cpu_irq_0_s0_writedata),              //                               .writedata
		.fingerprint_0_avalon_master_writedata   (processor0_0_fingerprint_0_avalon_master_writedata),                 //    fingerprint_0_avalon_master.writedata
		.fingerprint_0_avalon_master_write       (processor0_0_fingerprint_0_avalon_master_write),                     //                               .write
		.fingerprint_0_avalon_master_readdata    (processor0_0_fingerprint_0_avalon_master_readdata),                  //                               .readdata
		.fingerprint_0_avalon_master_waitrequest (processor0_0_fingerprint_0_avalon_master_waitrequest),               //                               .waitrequest
		.fingerprint_0_avalon_master_read        (processor0_0_fingerprint_0_avalon_master_read),                      //                               .read
		.fingerprint_0_avalon_master_address     (processor0_0_fingerprint_0_avalon_master_address),                   //                               .address
		.dma_0_control_port_slave_address        (mm_interconnect_1_processor0_0_dma_0_control_port_slave_address),    //       dma_0_control_port_slave.address
		.dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor0_0_dma_0_control_port_slave_chipselect), //                               .chipselect
		.dma_0_control_port_slave_readdata       (mm_interconnect_1_processor0_0_dma_0_control_port_slave_readdata),   //                               .readdata
		.dma_0_control_port_slave_write_n        (~mm_interconnect_1_processor0_0_dma_0_control_port_slave_write),     //                               .write_n
		.dma_0_control_port_slave_writedata      (mm_interconnect_1_processor0_0_dma_0_control_port_slave_writedata),  //                               .writedata
		.dma_0_irq_irq                           (irq_mapper_receiver0_irq),                                           //                      dma_0_irq.irq
		.out_system_bridge_m0_waitrequest        (processor0_0_out_system_bridge_m0_waitrequest),                      //           out_system_bridge_m0.waitrequest
		.out_system_bridge_m0_readdata           (processor0_0_out_system_bridge_m0_readdata),                         //                               .readdata
		.out_system_bridge_m0_readdatavalid      (processor0_0_out_system_bridge_m0_readdatavalid),                    //                               .readdatavalid
		.out_system_bridge_m0_burstcount         (processor0_0_out_system_bridge_m0_burstcount),                       //                               .burstcount
		.out_system_bridge_m0_writedata          (processor0_0_out_system_bridge_m0_writedata),                        //                               .writedata
		.out_system_bridge_m0_address            (processor0_0_out_system_bridge_m0_address),                          //                               .address
		.out_system_bridge_m0_write              (processor0_0_out_system_bridge_m0_write),                            //                               .write
		.out_system_bridge_m0_read               (processor0_0_out_system_bridge_m0_read),                             //                               .read
		.out_system_bridge_m0_byteenable         (processor0_0_out_system_bridge_m0_byteenable),                       //                               .byteenable
		.out_system_bridge_m0_debugaccess        (processor0_0_out_system_bridge_m0_debugaccess),                      //                               .debugaccess
		.cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_address),   //      cpu_oflow_irq_0_avs_oflow.address
		.cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_write),     //                               .write
		.cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_writedata), //                               .writedata
		.cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_read),      //                               .read
		.cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_readdata)   //                               .readdata
	);

	nios_fprint_processorM_0 processorm_0 (
		.philosopher_clk_in_clk                (clk_clk),                                               //             philosopher_clk_in.clk
		.outgoing_master_waitrequest           (processorm_0_outgoing_master_waitrequest),              //                outgoing_master.waitrequest
		.outgoing_master_readdata              (processorm_0_outgoing_master_readdata),                 //                               .readdata
		.outgoing_master_readdatavalid         (processorm_0_outgoing_master_readdatavalid),            //                               .readdatavalid
		.outgoing_master_burstcount            (processorm_0_outgoing_master_burstcount),               //                               .burstcount
		.outgoing_master_writedata             (processorm_0_outgoing_master_writedata),                //                               .writedata
		.outgoing_master_address               (processorm_0_outgoing_master_address),                  //                               .address
		.outgoing_master_write                 (processorm_0_outgoing_master_write),                    //                               .write
		.outgoing_master_read                  (processorm_0_outgoing_master_read),                     //                               .read
		.outgoing_master_byteenable            (processorm_0_outgoing_master_byteenable),               //                               .byteenable
		.outgoing_master_debugaccess           (processorm_0_outgoing_master_debugaccess),              //                               .debugaccess
		.button_pio_external_connection_export (),                                                      // button_pio_external_connection.export
		.cpu0_jtag_debug_module_reset_reset    (),                                                      //   cpu0_jtag_debug_module_reset.reset
		.reset_reset_n                         (reset_reset_n),                                         //                          reset.reset_n
		.fprint_irq_0_irq_export               (cfpu_0_irq_export),                                     //               fprint_irq_0_irq.export
		.cpu_irq_0_s0_address                  (mm_interconnect_1_processorm_0_cpu_irq_0_s0_address),   //                   cpu_irq_0_s0.address
		.cpu_irq_0_s0_write                    (mm_interconnect_1_processorm_0_cpu_irq_0_s0_write),     //                               .write
		.cpu_irq_0_s0_writedata                (mm_interconnect_1_processorm_0_cpu_irq_0_s0_writedata), //                               .writedata
		.dma_0_irq_receiver_irq_irq            (processorm_0_dma_0_irq_receiver_irq_irq)                //         dma_0_irq_receiver_irq.irq
	);

	nios_fprint_processor2_0 processor2_0 (
		.philosopher_clk_in_clk                  (clk_clk),                                                            //             philosopher_clk_in.clk
		.button_pio_external_connection_export   (),                                                                   // button_pio_external_connection.export
		.cpu0_jtag_debug_module_reset_reset      (),                                                                   //   cpu0_jtag_debug_module_reset.reset
		.reset_reset_n                           (reset_reset_n),                                                      //                          reset.reset_n
		.cpu_irq_0_s0_address                    (mm_interconnect_1_processor2_0_cpu_irq_0_s0_address),                //                   cpu_irq_0_s0.address
		.cpu_irq_0_s0_write                      (mm_interconnect_1_processor2_0_cpu_irq_0_s0_write),                  //                               .write
		.cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor2_0_cpu_irq_0_s0_writedata),              //                               .writedata
		.fingerprint_0_avalon_master_writedata   (processor2_0_fingerprint_0_avalon_master_writedata),                 //    fingerprint_0_avalon_master.writedata
		.fingerprint_0_avalon_master_write       (processor2_0_fingerprint_0_avalon_master_write),                     //                               .write
		.fingerprint_0_avalon_master_readdata    (processor2_0_fingerprint_0_avalon_master_readdata),                  //                               .readdata
		.fingerprint_0_avalon_master_waitrequest (processor2_0_fingerprint_0_avalon_master_waitrequest),               //                               .waitrequest
		.fingerprint_0_avalon_master_read        (processor2_0_fingerprint_0_avalon_master_read),                      //                               .read
		.fingerprint_0_avalon_master_address     (processor2_0_fingerprint_0_avalon_master_address),                   //                               .address
		.dma_0_control_port_slave_address        (mm_interconnect_1_processor2_0_dma_0_control_port_slave_address),    //       dma_0_control_port_slave.address
		.dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor2_0_dma_0_control_port_slave_chipselect), //                               .chipselect
		.dma_0_control_port_slave_readdata       (mm_interconnect_1_processor2_0_dma_0_control_port_slave_readdata),   //                               .readdata
		.dma_0_control_port_slave_write_n        (~mm_interconnect_1_processor2_0_dma_0_control_port_slave_write),     //                               .write_n
		.dma_0_control_port_slave_writedata      (mm_interconnect_1_processor2_0_dma_0_control_port_slave_writedata),  //                               .writedata
		.dma_0_irq_irq                           (irq_mapper_receiver2_irq),                                           //                      dma_0_irq.irq
		.out_system_bridge_m0_waitrequest        (processor2_0_out_system_bridge_m0_waitrequest),                      //           out_system_bridge_m0.waitrequest
		.out_system_bridge_m0_readdata           (processor2_0_out_system_bridge_m0_readdata),                         //                               .readdata
		.out_system_bridge_m0_readdatavalid      (processor2_0_out_system_bridge_m0_readdatavalid),                    //                               .readdatavalid
		.out_system_bridge_m0_burstcount         (processor2_0_out_system_bridge_m0_burstcount),                       //                               .burstcount
		.out_system_bridge_m0_writedata          (processor2_0_out_system_bridge_m0_writedata),                        //                               .writedata
		.out_system_bridge_m0_address            (processor2_0_out_system_bridge_m0_address),                          //                               .address
		.out_system_bridge_m0_write              (processor2_0_out_system_bridge_m0_write),                            //                               .write
		.out_system_bridge_m0_read               (processor2_0_out_system_bridge_m0_read),                             //                               .read
		.out_system_bridge_m0_byteenable         (processor2_0_out_system_bridge_m0_byteenable),                       //                               .byteenable
		.out_system_bridge_m0_debugaccess        (processor2_0_out_system_bridge_m0_debugaccess),                      //                               .debugaccess
		.cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_address),   //      cpu_oflow_irq_0_avs_oflow.address
		.cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_write),     //                               .write
		.cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_writedata), //                               .writedata
		.cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_read),      //                               .read
		.cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_readdata)   //                               .readdata
	);

	nios_fprint_processor3_0 processor3_0 (
		.philosopher_clk_in_clk                  (clk_clk),                                                            //             philosopher_clk_in.clk
		.button_pio_external_connection_export   (),                                                                   // button_pio_external_connection.export
		.cpu0_jtag_debug_module_reset_reset      (),                                                                   //   cpu0_jtag_debug_module_reset.reset
		.reset_reset_n                           (reset_reset_n),                                                      //                          reset.reset_n
		.cpu_irq_0_s0_address                    (mm_interconnect_1_processor3_0_cpu_irq_0_s0_address),                //                   cpu_irq_0_s0.address
		.cpu_irq_0_s0_write                      (mm_interconnect_1_processor3_0_cpu_irq_0_s0_write),                  //                               .write
		.cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor3_0_cpu_irq_0_s0_writedata),              //                               .writedata
		.fingerprint_0_avalon_master_writedata   (processor3_0_fingerprint_0_avalon_master_writedata),                 //    fingerprint_0_avalon_master.writedata
		.fingerprint_0_avalon_master_write       (processor3_0_fingerprint_0_avalon_master_write),                     //                               .write
		.fingerprint_0_avalon_master_readdata    (processor3_0_fingerprint_0_avalon_master_readdata),                  //                               .readdata
		.fingerprint_0_avalon_master_waitrequest (processor3_0_fingerprint_0_avalon_master_waitrequest),               //                               .waitrequest
		.fingerprint_0_avalon_master_read        (processor3_0_fingerprint_0_avalon_master_read),                      //                               .read
		.fingerprint_0_avalon_master_address     (processor3_0_fingerprint_0_avalon_master_address),                   //                               .address
		.dma_0_control_port_slave_address        (mm_interconnect_1_processor3_0_dma_0_control_port_slave_address),    //       dma_0_control_port_slave.address
		.dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor3_0_dma_0_control_port_slave_chipselect), //                               .chipselect
		.dma_0_control_port_slave_readdata       (mm_interconnect_1_processor3_0_dma_0_control_port_slave_readdata),   //                               .readdata
		.dma_0_control_port_slave_write_n        (~mm_interconnect_1_processor3_0_dma_0_control_port_slave_write),     //                               .write_n
		.dma_0_control_port_slave_writedata      (mm_interconnect_1_processor3_0_dma_0_control_port_slave_writedata),  //                               .writedata
		.dma_0_irq_irq                           (irq_mapper_receiver3_irq),                                           //                      dma_0_irq.irq
		.out_system_bridge_m0_waitrequest        (processor3_0_out_system_bridge_m0_waitrequest),                      //           out_system_bridge_m0.waitrequest
		.out_system_bridge_m0_readdata           (processor3_0_out_system_bridge_m0_readdata),                         //                               .readdata
		.out_system_bridge_m0_readdatavalid      (processor3_0_out_system_bridge_m0_readdatavalid),                    //                               .readdatavalid
		.out_system_bridge_m0_burstcount         (processor3_0_out_system_bridge_m0_burstcount),                       //                               .burstcount
		.out_system_bridge_m0_writedata          (processor3_0_out_system_bridge_m0_writedata),                        //                               .writedata
		.out_system_bridge_m0_address            (processor3_0_out_system_bridge_m0_address),                          //                               .address
		.out_system_bridge_m0_write              (processor3_0_out_system_bridge_m0_write),                            //                               .write
		.out_system_bridge_m0_read               (processor3_0_out_system_bridge_m0_read),                             //                               .read
		.out_system_bridge_m0_byteenable         (processor3_0_out_system_bridge_m0_byteenable),                       //                               .byteenable
		.out_system_bridge_m0_debugaccess        (processor3_0_out_system_bridge_m0_debugaccess),                      //                               .debugaccess
		.cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_address),   //      cpu_oflow_irq_0_avs_oflow.address
		.cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_write),     //                               .write
		.cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_writedata), //                               .writedata
		.cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_read),      //                               .read
		.cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_readdata)   //                               .readdata
	);

	nios_fprint_processor4_0 processor4_0 (
		.philosopher_clk_in_clk                  (clk_clk),                                                            //             philosopher_clk_in.clk
		.button_pio_external_connection_export   (),                                                                   // button_pio_external_connection.export
		.cpu0_jtag_debug_module_reset_reset      (),                                                                   //   cpu0_jtag_debug_module_reset.reset
		.reset_reset_n                           (reset_reset_n),                                                      //                          reset.reset_n
		.cpu_irq_0_s0_address                    (mm_interconnect_1_processor4_0_cpu_irq_0_s0_address),                //                   cpu_irq_0_s0.address
		.cpu_irq_0_s0_write                      (mm_interconnect_1_processor4_0_cpu_irq_0_s0_write),                  //                               .write
		.cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor4_0_cpu_irq_0_s0_writedata),              //                               .writedata
		.fingerprint_0_avalon_master_writedata   (processor4_0_fingerprint_0_avalon_master_writedata),                 //    fingerprint_0_avalon_master.writedata
		.fingerprint_0_avalon_master_write       (processor4_0_fingerprint_0_avalon_master_write),                     //                               .write
		.fingerprint_0_avalon_master_readdata    (processor4_0_fingerprint_0_avalon_master_readdata),                  //                               .readdata
		.fingerprint_0_avalon_master_waitrequest (processor4_0_fingerprint_0_avalon_master_waitrequest),               //                               .waitrequest
		.fingerprint_0_avalon_master_read        (processor4_0_fingerprint_0_avalon_master_read),                      //                               .read
		.fingerprint_0_avalon_master_address     (processor4_0_fingerprint_0_avalon_master_address),                   //                               .address
		.dma_0_control_port_slave_address        (mm_interconnect_1_processor4_0_dma_0_control_port_slave_address),    //       dma_0_control_port_slave.address
		.dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor4_0_dma_0_control_port_slave_chipselect), //                               .chipselect
		.dma_0_control_port_slave_readdata       (mm_interconnect_1_processor4_0_dma_0_control_port_slave_readdata),   //                               .readdata
		.dma_0_control_port_slave_write_n        (~mm_interconnect_1_processor4_0_dma_0_control_port_slave_write),     //                               .write_n
		.dma_0_control_port_slave_writedata      (mm_interconnect_1_processor4_0_dma_0_control_port_slave_writedata),  //                               .writedata
		.dma_0_irq_irq                           (irq_mapper_receiver4_irq),                                           //                      dma_0_irq.irq
		.out_system_bridge_m0_waitrequest        (processor4_0_out_system_bridge_m0_waitrequest),                      //           out_system_bridge_m0.waitrequest
		.out_system_bridge_m0_readdata           (processor4_0_out_system_bridge_m0_readdata),                         //                               .readdata
		.out_system_bridge_m0_readdatavalid      (processor4_0_out_system_bridge_m0_readdatavalid),                    //                               .readdatavalid
		.out_system_bridge_m0_burstcount         (processor4_0_out_system_bridge_m0_burstcount),                       //                               .burstcount
		.out_system_bridge_m0_writedata          (processor4_0_out_system_bridge_m0_writedata),                        //                               .writedata
		.out_system_bridge_m0_address            (processor4_0_out_system_bridge_m0_address),                          //                               .address
		.out_system_bridge_m0_write              (processor4_0_out_system_bridge_m0_write),                            //                               .write
		.out_system_bridge_m0_read               (processor4_0_out_system_bridge_m0_read),                             //                               .read
		.out_system_bridge_m0_byteenable         (processor4_0_out_system_bridge_m0_byteenable),                       //                               .byteenable
		.out_system_bridge_m0_debugaccess        (processor4_0_out_system_bridge_m0_debugaccess),                      //                               .debugaccess
		.cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_address),   //      cpu_oflow_irq_0_avs_oflow.address
		.cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_write),     //                               .write
		.cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_writedata), //                               .writedata
		.cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_read),      //                               .read
		.cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_readdata)   //                               .readdata
	);

	nios_fprint_processor5_0 processor5_0 (
		.philosopher_clk_in_clk                  (clk_clk),                                                            //             philosopher_clk_in.clk
		.button_pio_external_connection_export   (),                                                                   // button_pio_external_connection.export
		.cpu0_jtag_debug_module_reset_reset      (),                                                                   //   cpu0_jtag_debug_module_reset.reset
		.reset_reset_n                           (reset_reset_n),                                                      //                          reset.reset_n
		.cpu_irq_0_s0_address                    (mm_interconnect_1_processor5_0_cpu_irq_0_s0_address),                //                   cpu_irq_0_s0.address
		.cpu_irq_0_s0_write                      (mm_interconnect_1_processor5_0_cpu_irq_0_s0_write),                  //                               .write
		.cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor5_0_cpu_irq_0_s0_writedata),              //                               .writedata
		.fingerprint_0_avalon_master_writedata   (processor5_0_fingerprint_0_avalon_master_writedata),                 //    fingerprint_0_avalon_master.writedata
		.fingerprint_0_avalon_master_write       (processor5_0_fingerprint_0_avalon_master_write),                     //                               .write
		.fingerprint_0_avalon_master_readdata    (processor5_0_fingerprint_0_avalon_master_readdata),                  //                               .readdata
		.fingerprint_0_avalon_master_waitrequest (processor5_0_fingerprint_0_avalon_master_waitrequest),               //                               .waitrequest
		.fingerprint_0_avalon_master_read        (processor5_0_fingerprint_0_avalon_master_read),                      //                               .read
		.fingerprint_0_avalon_master_address     (processor5_0_fingerprint_0_avalon_master_address),                   //                               .address
		.dma_0_control_port_slave_address        (mm_interconnect_1_processor5_0_dma_0_control_port_slave_address),    //       dma_0_control_port_slave.address
		.dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor5_0_dma_0_control_port_slave_chipselect), //                               .chipselect
		.dma_0_control_port_slave_readdata       (mm_interconnect_1_processor5_0_dma_0_control_port_slave_readdata),   //                               .readdata
		.dma_0_control_port_slave_write_n        (~mm_interconnect_1_processor5_0_dma_0_control_port_slave_write),     //                               .write_n
		.dma_0_control_port_slave_writedata      (mm_interconnect_1_processor5_0_dma_0_control_port_slave_writedata),  //                               .writedata
		.dma_0_irq_irq                           (irq_mapper_receiver5_irq),                                           //                      dma_0_irq.irq
		.out_system_bridge_m0_waitrequest        (processor5_0_out_system_bridge_m0_waitrequest),                      //           out_system_bridge_m0.waitrequest
		.out_system_bridge_m0_readdata           (processor5_0_out_system_bridge_m0_readdata),                         //                               .readdata
		.out_system_bridge_m0_readdatavalid      (processor5_0_out_system_bridge_m0_readdatavalid),                    //                               .readdatavalid
		.out_system_bridge_m0_burstcount         (processor5_0_out_system_bridge_m0_burstcount),                       //                               .burstcount
		.out_system_bridge_m0_writedata          (processor5_0_out_system_bridge_m0_writedata),                        //                               .writedata
		.out_system_bridge_m0_address            (processor5_0_out_system_bridge_m0_address),                          //                               .address
		.out_system_bridge_m0_write              (processor5_0_out_system_bridge_m0_write),                            //                               .write
		.out_system_bridge_m0_read               (processor5_0_out_system_bridge_m0_read),                             //                               .read
		.out_system_bridge_m0_byteenable         (processor5_0_out_system_bridge_m0_byteenable),                       //                               .byteenable
		.out_system_bridge_m0_debugaccess        (processor5_0_out_system_bridge_m0_debugaccess),                      //                               .debugaccess
		.cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_address),   //      cpu_oflow_irq_0_avs_oflow.address
		.cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_write),     //                               .write
		.cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_writedata), //                               .writedata
		.cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_read),      //                               .read
		.cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_readdata)   //                               .readdata
	);

	nios_fprint_processor6_0 processor6_0 (
		.philosopher_clk_in_clk                  (clk_clk),                                                            //             philosopher_clk_in.clk
		.button_pio_external_connection_export   (),                                                                   // button_pio_external_connection.export
		.cpu0_jtag_debug_module_reset_reset      (),                                                                   //   cpu0_jtag_debug_module_reset.reset
		.reset_reset_n                           (reset_reset_n),                                                      //                          reset.reset_n
		.cpu_irq_0_s0_address                    (mm_interconnect_1_processor6_0_cpu_irq_0_s0_address),                //                   cpu_irq_0_s0.address
		.cpu_irq_0_s0_write                      (mm_interconnect_1_processor6_0_cpu_irq_0_s0_write),                  //                               .write
		.cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor6_0_cpu_irq_0_s0_writedata),              //                               .writedata
		.fingerprint_0_avalon_master_writedata   (processor6_0_fingerprint_0_avalon_master_writedata),                 //    fingerprint_0_avalon_master.writedata
		.fingerprint_0_avalon_master_write       (processor6_0_fingerprint_0_avalon_master_write),                     //                               .write
		.fingerprint_0_avalon_master_readdata    (processor6_0_fingerprint_0_avalon_master_readdata),                  //                               .readdata
		.fingerprint_0_avalon_master_waitrequest (processor6_0_fingerprint_0_avalon_master_waitrequest),               //                               .waitrequest
		.fingerprint_0_avalon_master_read        (processor6_0_fingerprint_0_avalon_master_read),                      //                               .read
		.fingerprint_0_avalon_master_address     (processor6_0_fingerprint_0_avalon_master_address),                   //                               .address
		.dma_0_control_port_slave_address        (mm_interconnect_1_processor6_0_dma_0_control_port_slave_address),    //       dma_0_control_port_slave.address
		.dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor6_0_dma_0_control_port_slave_chipselect), //                               .chipselect
		.dma_0_control_port_slave_readdata       (mm_interconnect_1_processor6_0_dma_0_control_port_slave_readdata),   //                               .readdata
		.dma_0_control_port_slave_write_n        (~mm_interconnect_1_processor6_0_dma_0_control_port_slave_write),     //                               .write_n
		.dma_0_control_port_slave_writedata      (mm_interconnect_1_processor6_0_dma_0_control_port_slave_writedata),  //                               .writedata
		.dma_0_irq_irq                           (irq_mapper_receiver6_irq),                                           //                      dma_0_irq.irq
		.out_system_bridge_m0_waitrequest        (processor6_0_out_system_bridge_m0_waitrequest),                      //           out_system_bridge_m0.waitrequest
		.out_system_bridge_m0_readdata           (processor6_0_out_system_bridge_m0_readdata),                         //                               .readdata
		.out_system_bridge_m0_readdatavalid      (processor6_0_out_system_bridge_m0_readdatavalid),                    //                               .readdatavalid
		.out_system_bridge_m0_burstcount         (processor6_0_out_system_bridge_m0_burstcount),                       //                               .burstcount
		.out_system_bridge_m0_writedata          (processor6_0_out_system_bridge_m0_writedata),                        //                               .writedata
		.out_system_bridge_m0_address            (processor6_0_out_system_bridge_m0_address),                          //                               .address
		.out_system_bridge_m0_write              (processor6_0_out_system_bridge_m0_write),                            //                               .write
		.out_system_bridge_m0_read               (processor6_0_out_system_bridge_m0_read),                             //                               .read
		.out_system_bridge_m0_byteenable         (processor6_0_out_system_bridge_m0_byteenable),                       //                               .byteenable
		.out_system_bridge_m0_debugaccess        (processor6_0_out_system_bridge_m0_debugaccess),                      //                               .debugaccess
		.cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_address),   //      cpu_oflow_irq_0_avs_oflow.address
		.cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_write),     //                               .write
		.cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_writedata), //                               .writedata
		.cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_read),      //                               .read
		.cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_readdata)   //                               .readdata
	);

	nios_fprint_processor7_0 processor7_0 (
		.philosopher_clk_in_clk                  (clk_clk),                                                            //             philosopher_clk_in.clk
		.button_pio_external_connection_export   (),                                                                   // button_pio_external_connection.export
		.cpu0_jtag_debug_module_reset_reset      (),                                                                   //   cpu0_jtag_debug_module_reset.reset
		.reset_reset_n                           (reset_reset_n),                                                      //                          reset.reset_n
		.cpu_irq_0_s0_address                    (mm_interconnect_1_processor7_0_cpu_irq_0_s0_address),                //                   cpu_irq_0_s0.address
		.cpu_irq_0_s0_write                      (mm_interconnect_1_processor7_0_cpu_irq_0_s0_write),                  //                               .write
		.cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor7_0_cpu_irq_0_s0_writedata),              //                               .writedata
		.fingerprint_0_avalon_master_writedata   (processor7_0_fingerprint_0_avalon_master_writedata),                 //    fingerprint_0_avalon_master.writedata
		.fingerprint_0_avalon_master_write       (processor7_0_fingerprint_0_avalon_master_write),                     //                               .write
		.fingerprint_0_avalon_master_readdata    (processor7_0_fingerprint_0_avalon_master_readdata),                  //                               .readdata
		.fingerprint_0_avalon_master_waitrequest (processor7_0_fingerprint_0_avalon_master_waitrequest),               //                               .waitrequest
		.fingerprint_0_avalon_master_read        (processor7_0_fingerprint_0_avalon_master_read),                      //                               .read
		.fingerprint_0_avalon_master_address     (processor7_0_fingerprint_0_avalon_master_address),                   //                               .address
		.dma_0_control_port_slave_address        (mm_interconnect_1_processor7_0_dma_0_control_port_slave_address),    //       dma_0_control_port_slave.address
		.dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor7_0_dma_0_control_port_slave_chipselect), //                               .chipselect
		.dma_0_control_port_slave_readdata       (mm_interconnect_1_processor7_0_dma_0_control_port_slave_readdata),   //                               .readdata
		.dma_0_control_port_slave_write_n        (~mm_interconnect_1_processor7_0_dma_0_control_port_slave_write),     //                               .write_n
		.dma_0_control_port_slave_writedata      (mm_interconnect_1_processor7_0_dma_0_control_port_slave_writedata),  //                               .writedata
		.dma_0_irq_irq                           (irq_mapper_receiver7_irq),                                           //                      dma_0_irq.irq
		.out_system_bridge_m0_waitrequest        (processor7_0_out_system_bridge_m0_waitrequest),                      //           out_system_bridge_m0.waitrequest
		.out_system_bridge_m0_readdata           (processor7_0_out_system_bridge_m0_readdata),                         //                               .readdata
		.out_system_bridge_m0_readdatavalid      (processor7_0_out_system_bridge_m0_readdatavalid),                    //                               .readdatavalid
		.out_system_bridge_m0_burstcount         (processor7_0_out_system_bridge_m0_burstcount),                       //                               .burstcount
		.out_system_bridge_m0_writedata          (processor7_0_out_system_bridge_m0_writedata),                        //                               .writedata
		.out_system_bridge_m0_address            (processor7_0_out_system_bridge_m0_address),                          //                               .address
		.out_system_bridge_m0_write              (processor7_0_out_system_bridge_m0_write),                            //                               .write
		.out_system_bridge_m0_read               (processor7_0_out_system_bridge_m0_read),                             //                               .read
		.out_system_bridge_m0_byteenable         (processor7_0_out_system_bridge_m0_byteenable),                       //                               .byteenable
		.out_system_bridge_m0_debugaccess        (processor7_0_out_system_bridge_m0_debugaccess),                      //                               .debugaccess
		.cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_address),   //      cpu_oflow_irq_0_avs_oflow.address
		.cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_write),     //                               .write
		.cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_writedata), //                               .writedata
		.cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_read),      //                               .read
		.cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_readdata)   //                               .readdata
	);

	nios_fprint_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                 (clk_clk),                                                 //                               clk_0_clk.clk
		.memory_0_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                          //    memory_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                          // mm_bridge_0_reset_reset_bridge_in_reset.reset
		.mm_bridge_0_m0_address                        (mm_bridge_0_m0_address),                                  //                          mm_bridge_0_m0.address
		.mm_bridge_0_m0_waitrequest                    (mm_bridge_0_m0_waitrequest),                              //                                        .waitrequest
		.mm_bridge_0_m0_burstcount                     (mm_bridge_0_m0_burstcount),                               //                                        .burstcount
		.mm_bridge_0_m0_byteenable                     (mm_bridge_0_m0_byteenable),                               //                                        .byteenable
		.mm_bridge_0_m0_read                           (mm_bridge_0_m0_read),                                     //                                        .read
		.mm_bridge_0_m0_readdata                       (mm_bridge_0_m0_readdata),                                 //                                        .readdata
		.mm_bridge_0_m0_readdatavalid                  (mm_bridge_0_m0_readdatavalid),                            //                                        .readdatavalid
		.mm_bridge_0_m0_write                          (mm_bridge_0_m0_write),                                    //                                        .write
		.mm_bridge_0_m0_writedata                      (mm_bridge_0_m0_writedata),                                //                                        .writedata
		.mm_bridge_0_m0_debugaccess                    (mm_bridge_0_m0_debugaccess),                              //                                        .debugaccess
		.cfpu_0_fprint_address                         (mm_interconnect_0_cfpu_0_fprint_address),                 //                           cfpu_0_fprint.address
		.cfpu_0_fprint_write                           (mm_interconnect_0_cfpu_0_fprint_write),                   //                                        .write
		.cfpu_0_fprint_writedata                       (mm_interconnect_0_cfpu_0_fprint_writedata),               //                                        .writedata
		.cfpu_0_fprint_waitrequest                     (mm_interconnect_0_cfpu_0_fprint_waitrequest),             //                                        .waitrequest
		.memory_0_mm_bridge_0_s0_address               (mm_interconnect_0_memory_0_mm_bridge_0_s0_address),       //                 memory_0_mm_bridge_0_s0.address
		.memory_0_mm_bridge_0_s0_write                 (mm_interconnect_0_memory_0_mm_bridge_0_s0_write),         //                                        .write
		.memory_0_mm_bridge_0_s0_read                  (mm_interconnect_0_memory_0_mm_bridge_0_s0_read),          //                                        .read
		.memory_0_mm_bridge_0_s0_readdata              (mm_interconnect_0_memory_0_mm_bridge_0_s0_readdata),      //                                        .readdata
		.memory_0_mm_bridge_0_s0_writedata             (mm_interconnect_0_memory_0_mm_bridge_0_s0_writedata),     //                                        .writedata
		.memory_0_mm_bridge_0_s0_burstcount            (mm_interconnect_0_memory_0_mm_bridge_0_s0_burstcount),    //                                        .burstcount
		.memory_0_mm_bridge_0_s0_byteenable            (mm_interconnect_0_memory_0_mm_bridge_0_s0_byteenable),    //                                        .byteenable
		.memory_0_mm_bridge_0_s0_readdatavalid         (mm_interconnect_0_memory_0_mm_bridge_0_s0_readdatavalid), //                                        .readdatavalid
		.memory_0_mm_bridge_0_s0_waitrequest           (mm_interconnect_0_memory_0_mm_bridge_0_s0_waitrequest),   //                                        .waitrequest
		.memory_0_mm_bridge_0_s0_debugaccess           (mm_interconnect_0_memory_0_mm_bridge_0_s0_debugaccess),   //                                        .debugaccess
		.sys_id_control_slave_address                  (mm_interconnect_0_sys_id_control_slave_address),          //                    sys_id_control_slave.address
		.sys_id_control_slave_readdata                 (mm_interconnect_0_sys_id_control_slave_readdata)          //                                        .readdata
	);

	nios_fprint_mm_interconnect_1 mm_interconnect_1 (
		.clk_0_clk_clk                                        (clk_clk),                                                            //                                clk_0_clk.clk
		.cfpu_0_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                                     //       cfpu_0_reset_reset_bridge_in_reset.reset
		.processor1_0_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                     // processor1_0_reset_reset_bridge_in_reset.reset
		.cfpu_0_oflow_address                                 (cfpu_0_oflow_address),                                               //                             cfpu_0_oflow.address
		.cfpu_0_oflow_waitrequest                             (cfpu_0_oflow_waitrequest),                                           //                                         .waitrequest
		.cfpu_0_oflow_write                                   (cfpu_0_oflow_write),                                                 //                                         .write
		.cfpu_0_oflow_writedata                               (cfpu_0_oflow_writedata),                                             //                                         .writedata
		.processor0_0_fingerprint_0_avalon_master_address     (processor0_0_fingerprint_0_avalon_master_address),                   // processor0_0_fingerprint_0_avalon_master.address
		.processor0_0_fingerprint_0_avalon_master_waitrequest (processor0_0_fingerprint_0_avalon_master_waitrequest),               //                                         .waitrequest
		.processor0_0_fingerprint_0_avalon_master_read        (processor0_0_fingerprint_0_avalon_master_read),                      //                                         .read
		.processor0_0_fingerprint_0_avalon_master_readdata    (processor0_0_fingerprint_0_avalon_master_readdata),                  //                                         .readdata
		.processor0_0_fingerprint_0_avalon_master_write       (processor0_0_fingerprint_0_avalon_master_write),                     //                                         .write
		.processor0_0_fingerprint_0_avalon_master_writedata   (processor0_0_fingerprint_0_avalon_master_writedata),                 //                                         .writedata
		.processor0_0_out_system_bridge_m0_address            (processor0_0_out_system_bridge_m0_address),                          //        processor0_0_out_system_bridge_m0.address
		.processor0_0_out_system_bridge_m0_waitrequest        (processor0_0_out_system_bridge_m0_waitrequest),                      //                                         .waitrequest
		.processor0_0_out_system_bridge_m0_burstcount         (processor0_0_out_system_bridge_m0_burstcount),                       //                                         .burstcount
		.processor0_0_out_system_bridge_m0_byteenable         (processor0_0_out_system_bridge_m0_byteenable),                       //                                         .byteenable
		.processor0_0_out_system_bridge_m0_read               (processor0_0_out_system_bridge_m0_read),                             //                                         .read
		.processor0_0_out_system_bridge_m0_readdata           (processor0_0_out_system_bridge_m0_readdata),                         //                                         .readdata
		.processor0_0_out_system_bridge_m0_readdatavalid      (processor0_0_out_system_bridge_m0_readdatavalid),                    //                                         .readdatavalid
		.processor0_0_out_system_bridge_m0_write              (processor0_0_out_system_bridge_m0_write),                            //                                         .write
		.processor0_0_out_system_bridge_m0_writedata          (processor0_0_out_system_bridge_m0_writedata),                        //                                         .writedata
		.processor0_0_out_system_bridge_m0_debugaccess        (processor0_0_out_system_bridge_m0_debugaccess),                      //                                         .debugaccess
		.processor1_0_fingerprint_0_avalon_master_address     (processor1_0_fingerprint_0_avalon_master_address),                   // processor1_0_fingerprint_0_avalon_master.address
		.processor1_0_fingerprint_0_avalon_master_waitrequest (processor1_0_fingerprint_0_avalon_master_waitrequest),               //                                         .waitrequest
		.processor1_0_fingerprint_0_avalon_master_read        (processor1_0_fingerprint_0_avalon_master_read),                      //                                         .read
		.processor1_0_fingerprint_0_avalon_master_readdata    (processor1_0_fingerprint_0_avalon_master_readdata),                  //                                         .readdata
		.processor1_0_fingerprint_0_avalon_master_write       (processor1_0_fingerprint_0_avalon_master_write),                     //                                         .write
		.processor1_0_fingerprint_0_avalon_master_writedata   (processor1_0_fingerprint_0_avalon_master_writedata),                 //                                         .writedata
		.processor1_0_outgoing_master_address                 (processor1_0_outgoing_master_address),                               //             processor1_0_outgoing_master.address
		.processor1_0_outgoing_master_waitrequest             (processor1_0_outgoing_master_waitrequest),                           //                                         .waitrequest
		.processor1_0_outgoing_master_burstcount              (processor1_0_outgoing_master_burstcount),                            //                                         .burstcount
		.processor1_0_outgoing_master_byteenable              (processor1_0_outgoing_master_byteenable),                            //                                         .byteenable
		.processor1_0_outgoing_master_read                    (processor1_0_outgoing_master_read),                                  //                                         .read
		.processor1_0_outgoing_master_readdata                (processor1_0_outgoing_master_readdata),                              //                                         .readdata
		.processor1_0_outgoing_master_readdatavalid           (processor1_0_outgoing_master_readdatavalid),                         //                                         .readdatavalid
		.processor1_0_outgoing_master_write                   (processor1_0_outgoing_master_write),                                 //                                         .write
		.processor1_0_outgoing_master_writedata               (processor1_0_outgoing_master_writedata),                             //                                         .writedata
		.processor1_0_outgoing_master_debugaccess             (processor1_0_outgoing_master_debugaccess),                           //                                         .debugaccess
		.processor2_0_fingerprint_0_avalon_master_address     (processor2_0_fingerprint_0_avalon_master_address),                   // processor2_0_fingerprint_0_avalon_master.address
		.processor2_0_fingerprint_0_avalon_master_waitrequest (processor2_0_fingerprint_0_avalon_master_waitrequest),               //                                         .waitrequest
		.processor2_0_fingerprint_0_avalon_master_read        (processor2_0_fingerprint_0_avalon_master_read),                      //                                         .read
		.processor2_0_fingerprint_0_avalon_master_readdata    (processor2_0_fingerprint_0_avalon_master_readdata),                  //                                         .readdata
		.processor2_0_fingerprint_0_avalon_master_write       (processor2_0_fingerprint_0_avalon_master_write),                     //                                         .write
		.processor2_0_fingerprint_0_avalon_master_writedata   (processor2_0_fingerprint_0_avalon_master_writedata),                 //                                         .writedata
		.processor2_0_out_system_bridge_m0_address            (processor2_0_out_system_bridge_m0_address),                          //        processor2_0_out_system_bridge_m0.address
		.processor2_0_out_system_bridge_m0_waitrequest        (processor2_0_out_system_bridge_m0_waitrequest),                      //                                         .waitrequest
		.processor2_0_out_system_bridge_m0_burstcount         (processor2_0_out_system_bridge_m0_burstcount),                       //                                         .burstcount
		.processor2_0_out_system_bridge_m0_byteenable         (processor2_0_out_system_bridge_m0_byteenable),                       //                                         .byteenable
		.processor2_0_out_system_bridge_m0_read               (processor2_0_out_system_bridge_m0_read),                             //                                         .read
		.processor2_0_out_system_bridge_m0_readdata           (processor2_0_out_system_bridge_m0_readdata),                         //                                         .readdata
		.processor2_0_out_system_bridge_m0_readdatavalid      (processor2_0_out_system_bridge_m0_readdatavalid),                    //                                         .readdatavalid
		.processor2_0_out_system_bridge_m0_write              (processor2_0_out_system_bridge_m0_write),                            //                                         .write
		.processor2_0_out_system_bridge_m0_writedata          (processor2_0_out_system_bridge_m0_writedata),                        //                                         .writedata
		.processor2_0_out_system_bridge_m0_debugaccess        (processor2_0_out_system_bridge_m0_debugaccess),                      //                                         .debugaccess
		.processor3_0_fingerprint_0_avalon_master_address     (processor3_0_fingerprint_0_avalon_master_address),                   // processor3_0_fingerprint_0_avalon_master.address
		.processor3_0_fingerprint_0_avalon_master_waitrequest (processor3_0_fingerprint_0_avalon_master_waitrequest),               //                                         .waitrequest
		.processor3_0_fingerprint_0_avalon_master_read        (processor3_0_fingerprint_0_avalon_master_read),                      //                                         .read
		.processor3_0_fingerprint_0_avalon_master_readdata    (processor3_0_fingerprint_0_avalon_master_readdata),                  //                                         .readdata
		.processor3_0_fingerprint_0_avalon_master_write       (processor3_0_fingerprint_0_avalon_master_write),                     //                                         .write
		.processor3_0_fingerprint_0_avalon_master_writedata   (processor3_0_fingerprint_0_avalon_master_writedata),                 //                                         .writedata
		.processor3_0_out_system_bridge_m0_address            (processor3_0_out_system_bridge_m0_address),                          //        processor3_0_out_system_bridge_m0.address
		.processor3_0_out_system_bridge_m0_waitrequest        (processor3_0_out_system_bridge_m0_waitrequest),                      //                                         .waitrequest
		.processor3_0_out_system_bridge_m0_burstcount         (processor3_0_out_system_bridge_m0_burstcount),                       //                                         .burstcount
		.processor3_0_out_system_bridge_m0_byteenable         (processor3_0_out_system_bridge_m0_byteenable),                       //                                         .byteenable
		.processor3_0_out_system_bridge_m0_read               (processor3_0_out_system_bridge_m0_read),                             //                                         .read
		.processor3_0_out_system_bridge_m0_readdata           (processor3_0_out_system_bridge_m0_readdata),                         //                                         .readdata
		.processor3_0_out_system_bridge_m0_readdatavalid      (processor3_0_out_system_bridge_m0_readdatavalid),                    //                                         .readdatavalid
		.processor3_0_out_system_bridge_m0_write              (processor3_0_out_system_bridge_m0_write),                            //                                         .write
		.processor3_0_out_system_bridge_m0_writedata          (processor3_0_out_system_bridge_m0_writedata),                        //                                         .writedata
		.processor3_0_out_system_bridge_m0_debugaccess        (processor3_0_out_system_bridge_m0_debugaccess),                      //                                         .debugaccess
		.processor4_0_fingerprint_0_avalon_master_address     (processor4_0_fingerprint_0_avalon_master_address),                   // processor4_0_fingerprint_0_avalon_master.address
		.processor4_0_fingerprint_0_avalon_master_waitrequest (processor4_0_fingerprint_0_avalon_master_waitrequest),               //                                         .waitrequest
		.processor4_0_fingerprint_0_avalon_master_read        (processor4_0_fingerprint_0_avalon_master_read),                      //                                         .read
		.processor4_0_fingerprint_0_avalon_master_readdata    (processor4_0_fingerprint_0_avalon_master_readdata),                  //                                         .readdata
		.processor4_0_fingerprint_0_avalon_master_write       (processor4_0_fingerprint_0_avalon_master_write),                     //                                         .write
		.processor4_0_fingerprint_0_avalon_master_writedata   (processor4_0_fingerprint_0_avalon_master_writedata),                 //                                         .writedata
		.processor4_0_out_system_bridge_m0_address            (processor4_0_out_system_bridge_m0_address),                          //        processor4_0_out_system_bridge_m0.address
		.processor4_0_out_system_bridge_m0_waitrequest        (processor4_0_out_system_bridge_m0_waitrequest),                      //                                         .waitrequest
		.processor4_0_out_system_bridge_m0_burstcount         (processor4_0_out_system_bridge_m0_burstcount),                       //                                         .burstcount
		.processor4_0_out_system_bridge_m0_byteenable         (processor4_0_out_system_bridge_m0_byteenable),                       //                                         .byteenable
		.processor4_0_out_system_bridge_m0_read               (processor4_0_out_system_bridge_m0_read),                             //                                         .read
		.processor4_0_out_system_bridge_m0_readdata           (processor4_0_out_system_bridge_m0_readdata),                         //                                         .readdata
		.processor4_0_out_system_bridge_m0_readdatavalid      (processor4_0_out_system_bridge_m0_readdatavalid),                    //                                         .readdatavalid
		.processor4_0_out_system_bridge_m0_write              (processor4_0_out_system_bridge_m0_write),                            //                                         .write
		.processor4_0_out_system_bridge_m0_writedata          (processor4_0_out_system_bridge_m0_writedata),                        //                                         .writedata
		.processor4_0_out_system_bridge_m0_debugaccess        (processor4_0_out_system_bridge_m0_debugaccess),                      //                                         .debugaccess
		.processor5_0_fingerprint_0_avalon_master_address     (processor5_0_fingerprint_0_avalon_master_address),                   // processor5_0_fingerprint_0_avalon_master.address
		.processor5_0_fingerprint_0_avalon_master_waitrequest (processor5_0_fingerprint_0_avalon_master_waitrequest),               //                                         .waitrequest
		.processor5_0_fingerprint_0_avalon_master_read        (processor5_0_fingerprint_0_avalon_master_read),                      //                                         .read
		.processor5_0_fingerprint_0_avalon_master_readdata    (processor5_0_fingerprint_0_avalon_master_readdata),                  //                                         .readdata
		.processor5_0_fingerprint_0_avalon_master_write       (processor5_0_fingerprint_0_avalon_master_write),                     //                                         .write
		.processor5_0_fingerprint_0_avalon_master_writedata   (processor5_0_fingerprint_0_avalon_master_writedata),                 //                                         .writedata
		.processor5_0_out_system_bridge_m0_address            (processor5_0_out_system_bridge_m0_address),                          //        processor5_0_out_system_bridge_m0.address
		.processor5_0_out_system_bridge_m0_waitrequest        (processor5_0_out_system_bridge_m0_waitrequest),                      //                                         .waitrequest
		.processor5_0_out_system_bridge_m0_burstcount         (processor5_0_out_system_bridge_m0_burstcount),                       //                                         .burstcount
		.processor5_0_out_system_bridge_m0_byteenable         (processor5_0_out_system_bridge_m0_byteenable),                       //                                         .byteenable
		.processor5_0_out_system_bridge_m0_read               (processor5_0_out_system_bridge_m0_read),                             //                                         .read
		.processor5_0_out_system_bridge_m0_readdata           (processor5_0_out_system_bridge_m0_readdata),                         //                                         .readdata
		.processor5_0_out_system_bridge_m0_readdatavalid      (processor5_0_out_system_bridge_m0_readdatavalid),                    //                                         .readdatavalid
		.processor5_0_out_system_bridge_m0_write              (processor5_0_out_system_bridge_m0_write),                            //                                         .write
		.processor5_0_out_system_bridge_m0_writedata          (processor5_0_out_system_bridge_m0_writedata),                        //                                         .writedata
		.processor5_0_out_system_bridge_m0_debugaccess        (processor5_0_out_system_bridge_m0_debugaccess),                      //                                         .debugaccess
		.processor6_0_fingerprint_0_avalon_master_address     (processor6_0_fingerprint_0_avalon_master_address),                   // processor6_0_fingerprint_0_avalon_master.address
		.processor6_0_fingerprint_0_avalon_master_waitrequest (processor6_0_fingerprint_0_avalon_master_waitrequest),               //                                         .waitrequest
		.processor6_0_fingerprint_0_avalon_master_read        (processor6_0_fingerprint_0_avalon_master_read),                      //                                         .read
		.processor6_0_fingerprint_0_avalon_master_readdata    (processor6_0_fingerprint_0_avalon_master_readdata),                  //                                         .readdata
		.processor6_0_fingerprint_0_avalon_master_write       (processor6_0_fingerprint_0_avalon_master_write),                     //                                         .write
		.processor6_0_fingerprint_0_avalon_master_writedata   (processor6_0_fingerprint_0_avalon_master_writedata),                 //                                         .writedata
		.processor6_0_out_system_bridge_m0_address            (processor6_0_out_system_bridge_m0_address),                          //        processor6_0_out_system_bridge_m0.address
		.processor6_0_out_system_bridge_m0_waitrequest        (processor6_0_out_system_bridge_m0_waitrequest),                      //                                         .waitrequest
		.processor6_0_out_system_bridge_m0_burstcount         (processor6_0_out_system_bridge_m0_burstcount),                       //                                         .burstcount
		.processor6_0_out_system_bridge_m0_byteenable         (processor6_0_out_system_bridge_m0_byteenable),                       //                                         .byteenable
		.processor6_0_out_system_bridge_m0_read               (processor6_0_out_system_bridge_m0_read),                             //                                         .read
		.processor6_0_out_system_bridge_m0_readdata           (processor6_0_out_system_bridge_m0_readdata),                         //                                         .readdata
		.processor6_0_out_system_bridge_m0_readdatavalid      (processor6_0_out_system_bridge_m0_readdatavalid),                    //                                         .readdatavalid
		.processor6_0_out_system_bridge_m0_write              (processor6_0_out_system_bridge_m0_write),                            //                                         .write
		.processor6_0_out_system_bridge_m0_writedata          (processor6_0_out_system_bridge_m0_writedata),                        //                                         .writedata
		.processor6_0_out_system_bridge_m0_debugaccess        (processor6_0_out_system_bridge_m0_debugaccess),                      //                                         .debugaccess
		.processor7_0_fingerprint_0_avalon_master_address     (processor7_0_fingerprint_0_avalon_master_address),                   // processor7_0_fingerprint_0_avalon_master.address
		.processor7_0_fingerprint_0_avalon_master_waitrequest (processor7_0_fingerprint_0_avalon_master_waitrequest),               //                                         .waitrequest
		.processor7_0_fingerprint_0_avalon_master_read        (processor7_0_fingerprint_0_avalon_master_read),                      //                                         .read
		.processor7_0_fingerprint_0_avalon_master_readdata    (processor7_0_fingerprint_0_avalon_master_readdata),                  //                                         .readdata
		.processor7_0_fingerprint_0_avalon_master_write       (processor7_0_fingerprint_0_avalon_master_write),                     //                                         .write
		.processor7_0_fingerprint_0_avalon_master_writedata   (processor7_0_fingerprint_0_avalon_master_writedata),                 //                                         .writedata
		.processor7_0_out_system_bridge_m0_address            (processor7_0_out_system_bridge_m0_address),                          //        processor7_0_out_system_bridge_m0.address
		.processor7_0_out_system_bridge_m0_waitrequest        (processor7_0_out_system_bridge_m0_waitrequest),                      //                                         .waitrequest
		.processor7_0_out_system_bridge_m0_burstcount         (processor7_0_out_system_bridge_m0_burstcount),                       //                                         .burstcount
		.processor7_0_out_system_bridge_m0_byteenable         (processor7_0_out_system_bridge_m0_byteenable),                       //                                         .byteenable
		.processor7_0_out_system_bridge_m0_read               (processor7_0_out_system_bridge_m0_read),                             //                                         .read
		.processor7_0_out_system_bridge_m0_readdata           (processor7_0_out_system_bridge_m0_readdata),                         //                                         .readdata
		.processor7_0_out_system_bridge_m0_readdatavalid      (processor7_0_out_system_bridge_m0_readdatavalid),                    //                                         .readdatavalid
		.processor7_0_out_system_bridge_m0_write              (processor7_0_out_system_bridge_m0_write),                            //                                         .write
		.processor7_0_out_system_bridge_m0_writedata          (processor7_0_out_system_bridge_m0_writedata),                        //                                         .writedata
		.processor7_0_out_system_bridge_m0_debugaccess        (processor7_0_out_system_bridge_m0_debugaccess),                      //                                         .debugaccess
		.processorM_0_outgoing_master_address                 (processorm_0_outgoing_master_address),                               //             processorM_0_outgoing_master.address
		.processorM_0_outgoing_master_waitrequest             (processorm_0_outgoing_master_waitrequest),                           //                                         .waitrequest
		.processorM_0_outgoing_master_burstcount              (processorm_0_outgoing_master_burstcount),                            //                                         .burstcount
		.processorM_0_outgoing_master_byteenable              (processorm_0_outgoing_master_byteenable),                            //                                         .byteenable
		.processorM_0_outgoing_master_read                    (processorm_0_outgoing_master_read),                                  //                                         .read
		.processorM_0_outgoing_master_readdata                (processorm_0_outgoing_master_readdata),                              //                                         .readdata
		.processorM_0_outgoing_master_readdatavalid           (processorm_0_outgoing_master_readdatavalid),                         //                                         .readdatavalid
		.processorM_0_outgoing_master_write                   (processorm_0_outgoing_master_write),                                 //                                         .write
		.processorM_0_outgoing_master_writedata               (processorm_0_outgoing_master_writedata),                             //                                         .writedata
		.processorM_0_outgoing_master_debugaccess             (processorm_0_outgoing_master_debugaccess),                           //                                         .debugaccess
		.cfpu_0_csr_address                                   (mm_interconnect_1_cfpu_0_csr_address),                               //                               cfpu_0_csr.address
		.cfpu_0_csr_write                                     (mm_interconnect_1_cfpu_0_csr_write),                                 //                                         .write
		.cfpu_0_csr_read                                      (mm_interconnect_1_cfpu_0_csr_read),                                  //                                         .read
		.cfpu_0_csr_readdata                                  (mm_interconnect_1_cfpu_0_csr_readdata),                              //                                         .readdata
		.cfpu_0_csr_writedata                                 (mm_interconnect_1_cfpu_0_csr_writedata),                             //                                         .writedata
		.cfpu_0_csr_waitrequest                               (mm_interconnect_1_cfpu_0_csr_waitrequest),                           //                                         .waitrequest
		.memory_0_memory_delay_0_csr_address                  (mm_interconnect_1_memory_0_memory_delay_0_csr_address),              //              memory_0_memory_delay_0_csr.address
		.memory_0_memory_delay_0_csr_write                    (mm_interconnect_1_memory_0_memory_delay_0_csr_write),                //                                         .write
		.memory_0_memory_delay_0_csr_writedata                (mm_interconnect_1_memory_0_memory_delay_0_csr_writedata),            //                                         .writedata
		.mm_bridge_0_s0_address                               (mm_interconnect_1_mm_bridge_0_s0_address),                           //                           mm_bridge_0_s0.address
		.mm_bridge_0_s0_write                                 (mm_interconnect_1_mm_bridge_0_s0_write),                             //                                         .write
		.mm_bridge_0_s0_read                                  (mm_interconnect_1_mm_bridge_0_s0_read),                              //                                         .read
		.mm_bridge_0_s0_readdata                              (mm_interconnect_1_mm_bridge_0_s0_readdata),                          //                                         .readdata
		.mm_bridge_0_s0_writedata                             (mm_interconnect_1_mm_bridge_0_s0_writedata),                         //                                         .writedata
		.mm_bridge_0_s0_burstcount                            (mm_interconnect_1_mm_bridge_0_s0_burstcount),                        //                                         .burstcount
		.mm_bridge_0_s0_byteenable                            (mm_interconnect_1_mm_bridge_0_s0_byteenable),                        //                                         .byteenable
		.mm_bridge_0_s0_readdatavalid                         (mm_interconnect_1_mm_bridge_0_s0_readdatavalid),                     //                                         .readdatavalid
		.mm_bridge_0_s0_waitrequest                           (mm_interconnect_1_mm_bridge_0_s0_waitrequest),                       //                                         .waitrequest
		.mm_bridge_0_s0_debugaccess                           (mm_interconnect_1_mm_bridge_0_s0_debugaccess),                       //                                         .debugaccess
		.mutex_0_s1_address                                   (mm_interconnect_1_mutex_0_s1_address),                               //                               mutex_0_s1.address
		.mutex_0_s1_write                                     (mm_interconnect_1_mutex_0_s1_write),                                 //                                         .write
		.mutex_0_s1_read                                      (mm_interconnect_1_mutex_0_s1_read),                                  //                                         .read
		.mutex_0_s1_readdata                                  (mm_interconnect_1_mutex_0_s1_readdata),                              //                                         .readdata
		.mutex_0_s1_writedata                                 (mm_interconnect_1_mutex_0_s1_writedata),                             //                                         .writedata
		.mutex_0_s1_chipselect                                (mm_interconnect_1_mutex_0_s1_chipselect),                            //                                         .chipselect
		.processor0_0_cpu_irq_0_s0_address                    (mm_interconnect_1_processor0_0_cpu_irq_0_s0_address),                //                processor0_0_cpu_irq_0_s0.address
		.processor0_0_cpu_irq_0_s0_write                      (mm_interconnect_1_processor0_0_cpu_irq_0_s0_write),                  //                                         .write
		.processor0_0_cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor0_0_cpu_irq_0_s0_writedata),              //                                         .writedata
		.processor0_0_cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_address),   //   processor0_0_cpu_oflow_irq_0_avs_oflow.address
		.processor0_0_cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_write),     //                                         .write
		.processor0_0_cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_read),      //                                         .read
		.processor0_0_cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_readdata),  //                                         .readdata
		.processor0_0_cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor0_0_cpu_oflow_irq_0_avs_oflow_writedata), //                                         .writedata
		.processor0_0_dma_0_control_port_slave_address        (mm_interconnect_1_processor0_0_dma_0_control_port_slave_address),    //    processor0_0_dma_0_control_port_slave.address
		.processor0_0_dma_0_control_port_slave_write          (mm_interconnect_1_processor0_0_dma_0_control_port_slave_write),      //                                         .write
		.processor0_0_dma_0_control_port_slave_readdata       (mm_interconnect_1_processor0_0_dma_0_control_port_slave_readdata),   //                                         .readdata
		.processor0_0_dma_0_control_port_slave_writedata      (mm_interconnect_1_processor0_0_dma_0_control_port_slave_writedata),  //                                         .writedata
		.processor0_0_dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor0_0_dma_0_control_port_slave_chipselect), //                                         .chipselect
		.processor1_0_cpu1_irq_0_s0_address                   (mm_interconnect_1_processor1_0_cpu1_irq_0_s0_address),               //               processor1_0_cpu1_irq_0_s0.address
		.processor1_0_cpu1_irq_0_s0_write                     (mm_interconnect_1_processor1_0_cpu1_irq_0_s0_write),                 //                                         .write
		.processor1_0_cpu1_irq_0_s0_writedata                 (mm_interconnect_1_processor1_0_cpu1_irq_0_s0_writedata),             //                                         .writedata
		.processor1_0_cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_address),   //   processor1_0_cpu_oflow_irq_0_avs_oflow.address
		.processor1_0_cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_write),     //                                         .write
		.processor1_0_cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_read),      //                                         .read
		.processor1_0_cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_readdata),  //                                         .readdata
		.processor1_0_cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor1_0_cpu_oflow_irq_0_avs_oflow_writedata), //                                         .writedata
		.processor1_0_dma_0_control_port_slave_address        (mm_interconnect_1_processor1_0_dma_0_control_port_slave_address),    //    processor1_0_dma_0_control_port_slave.address
		.processor1_0_dma_0_control_port_slave_write          (mm_interconnect_1_processor1_0_dma_0_control_port_slave_write),      //                                         .write
		.processor1_0_dma_0_control_port_slave_readdata       (mm_interconnect_1_processor1_0_dma_0_control_port_slave_readdata),   //                                         .readdata
		.processor1_0_dma_0_control_port_slave_writedata      (mm_interconnect_1_processor1_0_dma_0_control_port_slave_writedata),  //                                         .writedata
		.processor1_0_dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor1_0_dma_0_control_port_slave_chipselect), //                                         .chipselect
		.processor2_0_cpu_irq_0_s0_address                    (mm_interconnect_1_processor2_0_cpu_irq_0_s0_address),                //                processor2_0_cpu_irq_0_s0.address
		.processor2_0_cpu_irq_0_s0_write                      (mm_interconnect_1_processor2_0_cpu_irq_0_s0_write),                  //                                         .write
		.processor2_0_cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor2_0_cpu_irq_0_s0_writedata),              //                                         .writedata
		.processor2_0_cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_address),   //   processor2_0_cpu_oflow_irq_0_avs_oflow.address
		.processor2_0_cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_write),     //                                         .write
		.processor2_0_cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_read),      //                                         .read
		.processor2_0_cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_readdata),  //                                         .readdata
		.processor2_0_cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor2_0_cpu_oflow_irq_0_avs_oflow_writedata), //                                         .writedata
		.processor2_0_dma_0_control_port_slave_address        (mm_interconnect_1_processor2_0_dma_0_control_port_slave_address),    //    processor2_0_dma_0_control_port_slave.address
		.processor2_0_dma_0_control_port_slave_write          (mm_interconnect_1_processor2_0_dma_0_control_port_slave_write),      //                                         .write
		.processor2_0_dma_0_control_port_slave_readdata       (mm_interconnect_1_processor2_0_dma_0_control_port_slave_readdata),   //                                         .readdata
		.processor2_0_dma_0_control_port_slave_writedata      (mm_interconnect_1_processor2_0_dma_0_control_port_slave_writedata),  //                                         .writedata
		.processor2_0_dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor2_0_dma_0_control_port_slave_chipselect), //                                         .chipselect
		.processor3_0_cpu_irq_0_s0_address                    (mm_interconnect_1_processor3_0_cpu_irq_0_s0_address),                //                processor3_0_cpu_irq_0_s0.address
		.processor3_0_cpu_irq_0_s0_write                      (mm_interconnect_1_processor3_0_cpu_irq_0_s0_write),                  //                                         .write
		.processor3_0_cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor3_0_cpu_irq_0_s0_writedata),              //                                         .writedata
		.processor3_0_cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_address),   //   processor3_0_cpu_oflow_irq_0_avs_oflow.address
		.processor3_0_cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_write),     //                                         .write
		.processor3_0_cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_read),      //                                         .read
		.processor3_0_cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_readdata),  //                                         .readdata
		.processor3_0_cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor3_0_cpu_oflow_irq_0_avs_oflow_writedata), //                                         .writedata
		.processor3_0_dma_0_control_port_slave_address        (mm_interconnect_1_processor3_0_dma_0_control_port_slave_address),    //    processor3_0_dma_0_control_port_slave.address
		.processor3_0_dma_0_control_port_slave_write          (mm_interconnect_1_processor3_0_dma_0_control_port_slave_write),      //                                         .write
		.processor3_0_dma_0_control_port_slave_readdata       (mm_interconnect_1_processor3_0_dma_0_control_port_slave_readdata),   //                                         .readdata
		.processor3_0_dma_0_control_port_slave_writedata      (mm_interconnect_1_processor3_0_dma_0_control_port_slave_writedata),  //                                         .writedata
		.processor3_0_dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor3_0_dma_0_control_port_slave_chipselect), //                                         .chipselect
		.processor4_0_cpu_irq_0_s0_address                    (mm_interconnect_1_processor4_0_cpu_irq_0_s0_address),                //                processor4_0_cpu_irq_0_s0.address
		.processor4_0_cpu_irq_0_s0_write                      (mm_interconnect_1_processor4_0_cpu_irq_0_s0_write),                  //                                         .write
		.processor4_0_cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor4_0_cpu_irq_0_s0_writedata),              //                                         .writedata
		.processor4_0_cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_address),   //   processor4_0_cpu_oflow_irq_0_avs_oflow.address
		.processor4_0_cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_write),     //                                         .write
		.processor4_0_cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_read),      //                                         .read
		.processor4_0_cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_readdata),  //                                         .readdata
		.processor4_0_cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor4_0_cpu_oflow_irq_0_avs_oflow_writedata), //                                         .writedata
		.processor4_0_dma_0_control_port_slave_address        (mm_interconnect_1_processor4_0_dma_0_control_port_slave_address),    //    processor4_0_dma_0_control_port_slave.address
		.processor4_0_dma_0_control_port_slave_write          (mm_interconnect_1_processor4_0_dma_0_control_port_slave_write),      //                                         .write
		.processor4_0_dma_0_control_port_slave_readdata       (mm_interconnect_1_processor4_0_dma_0_control_port_slave_readdata),   //                                         .readdata
		.processor4_0_dma_0_control_port_slave_writedata      (mm_interconnect_1_processor4_0_dma_0_control_port_slave_writedata),  //                                         .writedata
		.processor4_0_dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor4_0_dma_0_control_port_slave_chipselect), //                                         .chipselect
		.processor5_0_cpu_irq_0_s0_address                    (mm_interconnect_1_processor5_0_cpu_irq_0_s0_address),                //                processor5_0_cpu_irq_0_s0.address
		.processor5_0_cpu_irq_0_s0_write                      (mm_interconnect_1_processor5_0_cpu_irq_0_s0_write),                  //                                         .write
		.processor5_0_cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor5_0_cpu_irq_0_s0_writedata),              //                                         .writedata
		.processor5_0_cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_address),   //   processor5_0_cpu_oflow_irq_0_avs_oflow.address
		.processor5_0_cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_write),     //                                         .write
		.processor5_0_cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_read),      //                                         .read
		.processor5_0_cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_readdata),  //                                         .readdata
		.processor5_0_cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor5_0_cpu_oflow_irq_0_avs_oflow_writedata), //                                         .writedata
		.processor5_0_dma_0_control_port_slave_address        (mm_interconnect_1_processor5_0_dma_0_control_port_slave_address),    //    processor5_0_dma_0_control_port_slave.address
		.processor5_0_dma_0_control_port_slave_write          (mm_interconnect_1_processor5_0_dma_0_control_port_slave_write),      //                                         .write
		.processor5_0_dma_0_control_port_slave_readdata       (mm_interconnect_1_processor5_0_dma_0_control_port_slave_readdata),   //                                         .readdata
		.processor5_0_dma_0_control_port_slave_writedata      (mm_interconnect_1_processor5_0_dma_0_control_port_slave_writedata),  //                                         .writedata
		.processor5_0_dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor5_0_dma_0_control_port_slave_chipselect), //                                         .chipselect
		.processor6_0_cpu_irq_0_s0_address                    (mm_interconnect_1_processor6_0_cpu_irq_0_s0_address),                //                processor6_0_cpu_irq_0_s0.address
		.processor6_0_cpu_irq_0_s0_write                      (mm_interconnect_1_processor6_0_cpu_irq_0_s0_write),                  //                                         .write
		.processor6_0_cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor6_0_cpu_irq_0_s0_writedata),              //                                         .writedata
		.processor6_0_cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_address),   //   processor6_0_cpu_oflow_irq_0_avs_oflow.address
		.processor6_0_cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_write),     //                                         .write
		.processor6_0_cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_read),      //                                         .read
		.processor6_0_cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_readdata),  //                                         .readdata
		.processor6_0_cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor6_0_cpu_oflow_irq_0_avs_oflow_writedata), //                                         .writedata
		.processor6_0_dma_0_control_port_slave_address        (mm_interconnect_1_processor6_0_dma_0_control_port_slave_address),    //    processor6_0_dma_0_control_port_slave.address
		.processor6_0_dma_0_control_port_slave_write          (mm_interconnect_1_processor6_0_dma_0_control_port_slave_write),      //                                         .write
		.processor6_0_dma_0_control_port_slave_readdata       (mm_interconnect_1_processor6_0_dma_0_control_port_slave_readdata),   //                                         .readdata
		.processor6_0_dma_0_control_port_slave_writedata      (mm_interconnect_1_processor6_0_dma_0_control_port_slave_writedata),  //                                         .writedata
		.processor6_0_dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor6_0_dma_0_control_port_slave_chipselect), //                                         .chipselect
		.processor7_0_cpu_irq_0_s0_address                    (mm_interconnect_1_processor7_0_cpu_irq_0_s0_address),                //                processor7_0_cpu_irq_0_s0.address
		.processor7_0_cpu_irq_0_s0_write                      (mm_interconnect_1_processor7_0_cpu_irq_0_s0_write),                  //                                         .write
		.processor7_0_cpu_irq_0_s0_writedata                  (mm_interconnect_1_processor7_0_cpu_irq_0_s0_writedata),              //                                         .writedata
		.processor7_0_cpu_oflow_irq_0_avs_oflow_address       (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_address),   //   processor7_0_cpu_oflow_irq_0_avs_oflow.address
		.processor7_0_cpu_oflow_irq_0_avs_oflow_write         (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_write),     //                                         .write
		.processor7_0_cpu_oflow_irq_0_avs_oflow_read          (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_read),      //                                         .read
		.processor7_0_cpu_oflow_irq_0_avs_oflow_readdata      (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_readdata),  //                                         .readdata
		.processor7_0_cpu_oflow_irq_0_avs_oflow_writedata     (mm_interconnect_1_processor7_0_cpu_oflow_irq_0_avs_oflow_writedata), //                                         .writedata
		.processor7_0_dma_0_control_port_slave_address        (mm_interconnect_1_processor7_0_dma_0_control_port_slave_address),    //    processor7_0_dma_0_control_port_slave.address
		.processor7_0_dma_0_control_port_slave_write          (mm_interconnect_1_processor7_0_dma_0_control_port_slave_write),      //                                         .write
		.processor7_0_dma_0_control_port_slave_readdata       (mm_interconnect_1_processor7_0_dma_0_control_port_slave_readdata),   //                                         .readdata
		.processor7_0_dma_0_control_port_slave_writedata      (mm_interconnect_1_processor7_0_dma_0_control_port_slave_writedata),  //                                         .writedata
		.processor7_0_dma_0_control_port_slave_chipselect     (mm_interconnect_1_processor7_0_dma_0_control_port_slave_chipselect), //                                         .chipselect
		.processorM_0_cpu_irq_0_s0_address                    (mm_interconnect_1_processorm_0_cpu_irq_0_s0_address),                //                processorM_0_cpu_irq_0_s0.address
		.processorM_0_cpu_irq_0_s0_write                      (mm_interconnect_1_processorm_0_cpu_irq_0_s0_write),                  //                                         .write
		.processorM_0_cpu_irq_0_s0_writedata                  (mm_interconnect_1_processorm_0_cpu_irq_0_s0_writedata),              //                                         .writedata
		.shared_memory_s1_address                             (mm_interconnect_1_shared_memory_s1_address),                         //                         shared_memory_s1.address
		.shared_memory_s1_write                               (mm_interconnect_1_shared_memory_s1_write),                           //                                         .write
		.shared_memory_s1_readdata                            (mm_interconnect_1_shared_memory_s1_readdata),                        //                                         .readdata
		.shared_memory_s1_writedata                           (mm_interconnect_1_shared_memory_s1_writedata),                       //                                         .writedata
		.shared_memory_s1_byteenable                          (mm_interconnect_1_shared_memory_s1_byteenable),                      //                                         .byteenable
		.shared_memory_s1_chipselect                          (mm_interconnect_1_shared_memory_s1_chipselect),                      //                                         .chipselect
		.shared_memory_s1_clken                               (mm_interconnect_1_shared_memory_s1_clken)                            //                                         .clken
	);

	nios_fprint_irq_mapper irq_mapper (
		.clk           (clk_clk),                                 //       clk.clk
		.reset         (rst_controller_reset_out_reset),          // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),                // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),                // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),                // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),                // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),                // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),                // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),                // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),                // receiver7.irq
		.sender_irq    (processorm_0_dma_0_irq_receiver_irq_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
