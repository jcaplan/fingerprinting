// nios_fprint_processorM_0.v

// Generated using ACDS version 13.1 162 at 2015.05.21.15:11:21

`timescale 1 ps / 1 ps
module nios_fprint_processorM_0 (
		input  wire        philosopher_clk_in_clk,                //             philosopher_clk_in.clk
		input  wire        outgoing_master_waitrequest,           //                outgoing_master.waitrequest
		input  wire [31:0] outgoing_master_readdata,              //                               .readdata
		input  wire        outgoing_master_readdatavalid,         //                               .readdatavalid
		output wire [0:0]  outgoing_master_burstcount,            //                               .burstcount
		output wire [31:0] outgoing_master_writedata,             //                               .writedata
		output wire [26:0] outgoing_master_address,               //                               .address
		output wire        outgoing_master_write,                 //                               .write
		output wire        outgoing_master_read,                  //                               .read
		output wire [3:0]  outgoing_master_byteenable,            //                               .byteenable
		output wire        outgoing_master_debugaccess,           //                               .debugaccess
		input  wire        button_pio_external_connection_export, // button_pio_external_connection.export
		output wire        cpu0_jtag_debug_module_reset_reset,    //   cpu0_jtag_debug_module_reset.reset
		input  wire        reset_reset_n,                         //                          reset.reset_n
		input  wire        fprint_irq_0_irq_export,               //               fprint_irq_0_irq.export
		input  wire [7:0]  cpu_irq_0_s0_address,                  //                   cpu_irq_0_s0.address
		input  wire        cpu_irq_0_s0_write,                    //                               .write
		input  wire [31:0] cpu_irq_0_s0_writedata,                //                               .writedata
		input  wire [0:0]  dma_0_irq_receiver_irq_irq,            //         dma_0_irq_receiver_irq.irq
		input  wire [0:0]  dma_1_irq_receiver_irq_irq             //         dma_1_irq_receiver_irq.irq
	);

	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_scratchpad_s1_writedata;                 // mm_interconnect_0:scratchpad_s1_writedata -> scratchpad:writedata
	wire  [11:0] mm_interconnect_0_scratchpad_s1_address;                   // mm_interconnect_0:scratchpad_s1_address -> scratchpad:address
	wire         mm_interconnect_0_scratchpad_s1_chipselect;                // mm_interconnect_0:scratchpad_s1_chipselect -> scratchpad:chipselect
	wire         mm_interconnect_0_scratchpad_s1_clken;                     // mm_interconnect_0:scratchpad_s1_clken -> scratchpad:clken
	wire         mm_interconnect_0_scratchpad_s1_write;                     // mm_interconnect_0:scratchpad_s1_write -> scratchpad:write
	wire  [31:0] mm_interconnect_0_scratchpad_s1_readdata;                  // scratchpad:readdata -> mm_interconnect_0:scratchpad_s1_readdata
	wire   [3:0] mm_interconnect_0_scratchpad_s1_byteenable;                // mm_interconnect_0:scratchpad_s1_byteenable -> scratchpad:byteenable
	wire         mm_interconnect_0_out_system_bridge_s0_waitrequest;        // out_system_bridge:s0_waitrequest -> mm_interconnect_0:out_system_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_out_system_bridge_s0_burstcount;         // mm_interconnect_0:out_system_bridge_s0_burstcount -> out_system_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_writedata;          // mm_interconnect_0:out_system_bridge_s0_writedata -> out_system_bridge:s0_writedata
	wire  [26:0] mm_interconnect_0_out_system_bridge_s0_address;            // mm_interconnect_0:out_system_bridge_s0_address -> out_system_bridge:s0_address
	wire         mm_interconnect_0_out_system_bridge_s0_write;              // mm_interconnect_0:out_system_bridge_s0_write -> out_system_bridge:s0_write
	wire         mm_interconnect_0_out_system_bridge_s0_read;               // mm_interconnect_0:out_system_bridge_s0_read -> out_system_bridge:s0_read
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_readdata;           // out_system_bridge:s0_readdata -> mm_interconnect_0:out_system_bridge_s0_readdata
	wire         mm_interconnect_0_out_system_bridge_s0_debugaccess;        // mm_interconnect_0:out_system_bridge_s0_debugaccess -> out_system_bridge:s0_debugaccess
	wire         mm_interconnect_0_out_system_bridge_s0_readdatavalid;      // out_system_bridge:s0_readdatavalid -> mm_interconnect_0:out_system_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_out_system_bridge_s0_byteenable;         // mm_interconnect_0:out_system_bridge_s0_byteenable -> out_system_bridge:s0_byteenable
	wire  [31:0] mm_interconnect_0_button_pio_s1_writedata;                 // mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	wire   [1:0] mm_interconnect_0_button_pio_s1_address;                   // mm_interconnect_0:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_0_button_pio_s1_chipselect;                // mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	wire         mm_interconnect_0_button_pio_s1_write;                     // mm_interconnect_0:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_0_button_pio_s1_readdata;                  // button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	wire         cpum_instruction_master_waitrequest;                       // mm_interconnect_0:cpuM_instruction_master_waitrequest -> cpuM:i_waitrequest
	wire  [27:0] cpum_instruction_master_address;                           // cpuM:i_address -> mm_interconnect_0:cpuM_instruction_master_address
	wire         cpum_instruction_master_read;                              // cpuM:i_read -> mm_interconnect_0:cpuM_instruction_master_read
	wire  [31:0] cpum_instruction_master_readdata;                          // mm_interconnect_0:cpuM_instruction_master_readdata -> cpuM:i_readdata
	wire         cpum_instruction_master_readdatavalid;                     // mm_interconnect_0:cpuM_instruction_master_readdatavalid -> cpuM:i_readdatavalid
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire         cpum_data_master_waitrequest;                              // mm_interconnect_0:cpuM_data_master_waitrequest -> cpuM:d_waitrequest
	wire  [31:0] cpum_data_master_writedata;                                // cpuM:d_writedata -> mm_interconnect_0:cpuM_data_master_writedata
	wire  [27:0] cpum_data_master_address;                                  // cpuM:d_address -> mm_interconnect_0:cpuM_data_master_address
	wire         cpum_data_master_write;                                    // cpuM:d_write -> mm_interconnect_0:cpuM_data_master_write
	wire         cpum_data_master_read;                                     // cpuM:d_read -> mm_interconnect_0:cpuM_data_master_read
	wire  [31:0] cpum_data_master_readdata;                                 // mm_interconnect_0:cpuM_data_master_readdata -> cpuM:d_readdata
	wire         cpum_data_master_debugaccess;                              // cpuM:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpuM_data_master_debugaccess
	wire   [3:0] cpum_data_master_byteenable;                               // cpuM:d_byteenable -> mm_interconnect_0:cpuM_data_master_byteenable
	wire         mm_interconnect_0_cpum_jtag_debug_module_waitrequest;      // cpuM:jtag_debug_module_waitrequest -> mm_interconnect_0:cpuM_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpum_jtag_debug_module_writedata;        // mm_interconnect_0:cpuM_jtag_debug_module_writedata -> cpuM:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpum_jtag_debug_module_address;          // mm_interconnect_0:cpuM_jtag_debug_module_address -> cpuM:jtag_debug_module_address
	wire         mm_interconnect_0_cpum_jtag_debug_module_write;            // mm_interconnect_0:cpuM_jtag_debug_module_write -> cpuM:jtag_debug_module_write
	wire         mm_interconnect_0_cpum_jtag_debug_module_read;             // mm_interconnect_0:cpuM_jtag_debug_module_read -> cpuM:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpum_jtag_debug_module_readdata;         // cpuM:jtag_debug_module_readdata -> mm_interconnect_0:cpuM_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpum_jtag_debug_module_debugaccess;      // mm_interconnect_0:cpuM_jtag_debug_module_debugaccess -> cpuM:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpum_jtag_debug_module_byteenable;       // mm_interconnect_0:cpuM_jtag_debug_module_byteenable -> cpuM:jtag_debug_module_byteenable
	wire  [15:0] mm_interconnect_0_timestamp_s1_writedata;                  // mm_interconnect_0:timestamp_s1_writedata -> timestamp:writedata
	wire   [3:0] mm_interconnect_0_timestamp_s1_address;                    // mm_interconnect_0:timestamp_s1_address -> timestamp:address
	wire         mm_interconnect_0_timestamp_s1_chipselect;                 // mm_interconnect_0:timestamp_s1_chipselect -> timestamp:chipselect
	wire         mm_interconnect_0_timestamp_s1_write;                      // mm_interconnect_0:timestamp_s1_write -> timestamp:write_n
	wire  [15:0] mm_interconnect_0_timestamp_s1_readdata;                   // timestamp:readdata -> mm_interconnect_0:timestamp_s1_readdata
	wire         irq_mapper_receiver0_irq;                                  // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // button_pio:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // cpu_irq_0:ins_irq0_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // fprint_irq_0:irq_out -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                  // dma_0_irq:sender0_irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                  // dma_1_irq:sender0_irq -> irq_mapper:receiver6_irq
	wire  [31:0] cpum_d_irq_irq;                                            // irq_mapper:sender_irq -> cpuM:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [button_pio:reset_n, cpuM:reset_n, cpu_irq_0:reset, dma_0_irq:reset, dma_1_irq:reset, fprint_irq_0:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpuM_reset_n_reset_bridge_in_reset_reset, out_system_bridge:reset, rst_translator:in_reset, scratchpad:reset, timer:reset_n, timestamp:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpuM:reset_req, rst_translator:reset_req_in, scratchpad:reset_req]

	nios_fprint_processorM_0_cpuM cpum (
		.clk                                   (philosopher_clk_in_clk),                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (cpum_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpum_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpum_data_master_read),                                //                          .read
		.d_readdata                            (cpum_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpum_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpum_data_master_write),                               //                          .write
		.d_writedata                           (cpum_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpum_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpum_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpum_instruction_master_read),                         //                          .read
		.i_readdata                            (cpum_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpum_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpum_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpum_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpum_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpum_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpum_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpum_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpum_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpum_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpum_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpum_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (27),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) out_system_bridge (
		.clk              (philosopher_clk_in_clk),                               //   clk.clk
		.reset            (rst_controller_reset_out_reset),                       // reset.reset
		.s0_waitrequest   (mm_interconnect_0_out_system_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_out_system_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_out_system_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_out_system_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_out_system_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_out_system_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_out_system_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_out_system_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_out_system_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_out_system_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (outgoing_master_waitrequest),                          //    m0.waitrequest
		.m0_readdata      (outgoing_master_readdata),                             //      .readdata
		.m0_readdatavalid (outgoing_master_readdatavalid),                        //      .readdatavalid
		.m0_burstcount    (outgoing_master_burstcount),                           //      .burstcount
		.m0_writedata     (outgoing_master_writedata),                            //      .writedata
		.m0_address       (outgoing_master_address),                              //      .address
		.m0_write         (outgoing_master_write),                                //      .write
		.m0_read          (outgoing_master_read),                                 //      .read
		.m0_byteenable    (outgoing_master_byteenable),                           //      .byteenable
		.m0_debugaccess   (outgoing_master_debugaccess)                           //      .debugaccess
	);

	nios_fprint_processor1_0_timer timer (
		.clk        (philosopher_clk_in_clk),                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	nios_fprint_processor1_0_jtag_uart jtag_uart (
		.clk            (philosopher_clk_in_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	nios_fprint_processor1_0_button_pio button_pio (
		.clk        (philosopher_clk_in_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                    //                 irq.irq
	);

	cpu_irq cpu_irq_0 (
		.avs_s0_address   (cpu_irq_0_s0_address),           //    s0.address
		.avs_s0_write     (cpu_irq_0_s0_write),             //      .write
		.avs_s0_writedata (cpu_irq_0_s0_writedata),         //      .writedata
		.clk              (philosopher_clk_in_clk),         // clock.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.ins_irq0_irq     (irq_mapper_receiver3_irq)        //  irq0.irq
	);

	nios_fprint_processor1_0_timestamp timestamp (
		.clk        (philosopher_clk_in_clk),                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_timestamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timestamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timestamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timestamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timestamp_s1_write),     //      .write_n
		.irq        ()                                           //   irq.irq
	);

	fprint_irq fprint_irq_0 (
		.irq_out (irq_mapper_receiver4_irq),       // interrupt_sender.irq
		.irq     (fprint_irq_0_irq_export),        //              irq.export
		.clk     (philosopher_clk_in_clk),         //            clock.clk
		.reset   (rst_controller_reset_out_reset)  //            reset.reset
	);

	altera_irq_bridge #(
		.IRQ_WIDTH (1)
	) dma_0_irq (
		.clk          (philosopher_clk_in_clk),         //          clk.clk
		.receiver_irq (dma_0_irq_receiver_irq_irq),     // receiver_irq.irq
		.reset        (rst_controller_reset_out_reset), //    clk_reset.reset
		.sender0_irq  (irq_mapper_receiver5_irq),       //  sender0_irq.irq
		.sender1_irq  (),                               //  (terminated)
		.sender2_irq  (),                               //  (terminated)
		.sender3_irq  (),                               //  (terminated)
		.sender4_irq  (),                               //  (terminated)
		.sender5_irq  (),                               //  (terminated)
		.sender6_irq  (),                               //  (terminated)
		.sender7_irq  (),                               //  (terminated)
		.sender8_irq  (),                               //  (terminated)
		.sender9_irq  (),                               //  (terminated)
		.sender10_irq (),                               //  (terminated)
		.sender11_irq (),                               //  (terminated)
		.sender12_irq (),                               //  (terminated)
		.sender13_irq (),                               //  (terminated)
		.sender14_irq (),                               //  (terminated)
		.sender15_irq (),                               //  (terminated)
		.sender16_irq (),                               //  (terminated)
		.sender17_irq (),                               //  (terminated)
		.sender18_irq (),                               //  (terminated)
		.sender19_irq (),                               //  (terminated)
		.sender20_irq (),                               //  (terminated)
		.sender21_irq (),                               //  (terminated)
		.sender22_irq (),                               //  (terminated)
		.sender23_irq (),                               //  (terminated)
		.sender24_irq (),                               //  (terminated)
		.sender25_irq (),                               //  (terminated)
		.sender26_irq (),                               //  (terminated)
		.sender27_irq (),                               //  (terminated)
		.sender28_irq (),                               //  (terminated)
		.sender29_irq (),                               //  (terminated)
		.sender30_irq (),                               //  (terminated)
		.sender31_irq ()                                //  (terminated)
	);

	altera_irq_bridge #(
		.IRQ_WIDTH (1)
	) dma_1_irq (
		.clk          (philosopher_clk_in_clk),         //          clk.clk
		.receiver_irq (dma_1_irq_receiver_irq_irq),     // receiver_irq.irq
		.reset        (rst_controller_reset_out_reset), //    clk_reset.reset
		.sender0_irq  (irq_mapper_receiver6_irq),       //  sender0_irq.irq
		.sender1_irq  (),                               //  (terminated)
		.sender2_irq  (),                               //  (terminated)
		.sender3_irq  (),                               //  (terminated)
		.sender4_irq  (),                               //  (terminated)
		.sender5_irq  (),                               //  (terminated)
		.sender6_irq  (),                               //  (terminated)
		.sender7_irq  (),                               //  (terminated)
		.sender8_irq  (),                               //  (terminated)
		.sender9_irq  (),                               //  (terminated)
		.sender10_irq (),                               //  (terminated)
		.sender11_irq (),                               //  (terminated)
		.sender12_irq (),                               //  (terminated)
		.sender13_irq (),                               //  (terminated)
		.sender14_irq (),                               //  (terminated)
		.sender15_irq (),                               //  (terminated)
		.sender16_irq (),                               //  (terminated)
		.sender17_irq (),                               //  (terminated)
		.sender18_irq (),                               //  (terminated)
		.sender19_irq (),                               //  (terminated)
		.sender20_irq (),                               //  (terminated)
		.sender21_irq (),                               //  (terminated)
		.sender22_irq (),                               //  (terminated)
		.sender23_irq (),                               //  (terminated)
		.sender24_irq (),                               //  (terminated)
		.sender25_irq (),                               //  (terminated)
		.sender26_irq (),                               //  (terminated)
		.sender27_irq (),                               //  (terminated)
		.sender28_irq (),                               //  (terminated)
		.sender29_irq (),                               //  (terminated)
		.sender30_irq (),                               //  (terminated)
		.sender31_irq ()                                //  (terminated)
	);

	nios_fprint_processorM_0_scratchpad scratchpad (
		.clk        (philosopher_clk_in_clk),                     //   clk1.clk
		.address    (mm_interconnect_0_scratchpad_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_scratchpad_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_scratchpad_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_scratchpad_s1_write),      //       .write
		.readdata   (mm_interconnect_0_scratchpad_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_scratchpad_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_scratchpad_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	nios_fprint_processorM_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                              (philosopher_clk_in_clk),                                    //                            clk_clk.clk
		.cpuM_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpuM_reset_n_reset_bridge_in_reset.reset
		.cpuM_data_master_address                 (cpum_data_master_address),                                  //                   cpuM_data_master.address
		.cpuM_data_master_waitrequest             (cpum_data_master_waitrequest),                              //                                   .waitrequest
		.cpuM_data_master_byteenable              (cpum_data_master_byteenable),                               //                                   .byteenable
		.cpuM_data_master_read                    (cpum_data_master_read),                                     //                                   .read
		.cpuM_data_master_readdata                (cpum_data_master_readdata),                                 //                                   .readdata
		.cpuM_data_master_write                   (cpum_data_master_write),                                    //                                   .write
		.cpuM_data_master_writedata               (cpum_data_master_writedata),                                //                                   .writedata
		.cpuM_data_master_debugaccess             (cpum_data_master_debugaccess),                              //                                   .debugaccess
		.cpuM_instruction_master_address          (cpum_instruction_master_address),                           //            cpuM_instruction_master.address
		.cpuM_instruction_master_waitrequest      (cpum_instruction_master_waitrequest),                       //                                   .waitrequest
		.cpuM_instruction_master_read             (cpum_instruction_master_read),                              //                                   .read
		.cpuM_instruction_master_readdata         (cpum_instruction_master_readdata),                          //                                   .readdata
		.cpuM_instruction_master_readdatavalid    (cpum_instruction_master_readdatavalid),                     //                                   .readdatavalid
		.button_pio_s1_address                    (mm_interconnect_0_button_pio_s1_address),                   //                      button_pio_s1.address
		.button_pio_s1_write                      (mm_interconnect_0_button_pio_s1_write),                     //                                   .write
		.button_pio_s1_readdata                   (mm_interconnect_0_button_pio_s1_readdata),                  //                                   .readdata
		.button_pio_s1_writedata                  (mm_interconnect_0_button_pio_s1_writedata),                 //                                   .writedata
		.button_pio_s1_chipselect                 (mm_interconnect_0_button_pio_s1_chipselect),                //                                   .chipselect
		.cpuM_jtag_debug_module_address           (mm_interconnect_0_cpum_jtag_debug_module_address),          //             cpuM_jtag_debug_module.address
		.cpuM_jtag_debug_module_write             (mm_interconnect_0_cpum_jtag_debug_module_write),            //                                   .write
		.cpuM_jtag_debug_module_read              (mm_interconnect_0_cpum_jtag_debug_module_read),             //                                   .read
		.cpuM_jtag_debug_module_readdata          (mm_interconnect_0_cpum_jtag_debug_module_readdata),         //                                   .readdata
		.cpuM_jtag_debug_module_writedata         (mm_interconnect_0_cpum_jtag_debug_module_writedata),        //                                   .writedata
		.cpuM_jtag_debug_module_byteenable        (mm_interconnect_0_cpum_jtag_debug_module_byteenable),       //                                   .byteenable
		.cpuM_jtag_debug_module_waitrequest       (mm_interconnect_0_cpum_jtag_debug_module_waitrequest),      //                                   .waitrequest
		.cpuM_jtag_debug_module_debugaccess       (mm_interconnect_0_cpum_jtag_debug_module_debugaccess),      //                                   .debugaccess
		.jtag_uart_avalon_jtag_slave_address      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                   .write
		.jtag_uart_avalon_jtag_slave_read         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                   .read
		.jtag_uart_avalon_jtag_slave_readdata     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.out_system_bridge_s0_address             (mm_interconnect_0_out_system_bridge_s0_address),            //               out_system_bridge_s0.address
		.out_system_bridge_s0_write               (mm_interconnect_0_out_system_bridge_s0_write),              //                                   .write
		.out_system_bridge_s0_read                (mm_interconnect_0_out_system_bridge_s0_read),               //                                   .read
		.out_system_bridge_s0_readdata            (mm_interconnect_0_out_system_bridge_s0_readdata),           //                                   .readdata
		.out_system_bridge_s0_writedata           (mm_interconnect_0_out_system_bridge_s0_writedata),          //                                   .writedata
		.out_system_bridge_s0_burstcount          (mm_interconnect_0_out_system_bridge_s0_burstcount),         //                                   .burstcount
		.out_system_bridge_s0_byteenable          (mm_interconnect_0_out_system_bridge_s0_byteenable),         //                                   .byteenable
		.out_system_bridge_s0_readdatavalid       (mm_interconnect_0_out_system_bridge_s0_readdatavalid),      //                                   .readdatavalid
		.out_system_bridge_s0_waitrequest         (mm_interconnect_0_out_system_bridge_s0_waitrequest),        //                                   .waitrequest
		.out_system_bridge_s0_debugaccess         (mm_interconnect_0_out_system_bridge_s0_debugaccess),        //                                   .debugaccess
		.scratchpad_s1_address                    (mm_interconnect_0_scratchpad_s1_address),                   //                      scratchpad_s1.address
		.scratchpad_s1_write                      (mm_interconnect_0_scratchpad_s1_write),                     //                                   .write
		.scratchpad_s1_readdata                   (mm_interconnect_0_scratchpad_s1_readdata),                  //                                   .readdata
		.scratchpad_s1_writedata                  (mm_interconnect_0_scratchpad_s1_writedata),                 //                                   .writedata
		.scratchpad_s1_byteenable                 (mm_interconnect_0_scratchpad_s1_byteenable),                //                                   .byteenable
		.scratchpad_s1_chipselect                 (mm_interconnect_0_scratchpad_s1_chipselect),                //                                   .chipselect
		.scratchpad_s1_clken                      (mm_interconnect_0_scratchpad_s1_clken),                     //                                   .clken
		.timer_s1_address                         (mm_interconnect_0_timer_s1_address),                        //                           timer_s1.address
		.timer_s1_write                           (mm_interconnect_0_timer_s1_write),                          //                                   .write
		.timer_s1_readdata                        (mm_interconnect_0_timer_s1_readdata),                       //                                   .readdata
		.timer_s1_writedata                       (mm_interconnect_0_timer_s1_writedata),                      //                                   .writedata
		.timer_s1_chipselect                      (mm_interconnect_0_timer_s1_chipselect),                     //                                   .chipselect
		.timestamp_s1_address                     (mm_interconnect_0_timestamp_s1_address),                    //                       timestamp_s1.address
		.timestamp_s1_write                       (mm_interconnect_0_timestamp_s1_write),                      //                                   .write
		.timestamp_s1_readdata                    (mm_interconnect_0_timestamp_s1_readdata),                   //                                   .readdata
		.timestamp_s1_writedata                   (mm_interconnect_0_timestamp_s1_writedata),                  //                                   .writedata
		.timestamp_s1_chipselect                  (mm_interconnect_0_timestamp_s1_chipselect)                  //                                   .chipselect
	);

	nios_fprint_processorM_0_irq_mapper irq_mapper (
		.clk           (philosopher_clk_in_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.sender_irq    (cpum_d_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (philosopher_clk_in_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
