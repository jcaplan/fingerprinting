library verilog;
use verilog.vl_types.all;
entity tb_oflow_registers is
end tb_oflow_registers;
