// nios_fprint_processorMonitor.v

// Generated using ACDS version 13.1 162 at 2014.07.12.16:57:40

`timescale 1 ps / 1 ps
module nios_fprint_processorMonitor (
		input  wire        philosopher_clk_in_clk,                //             philosopher_clk_in.clk
		input  wire        outgoing_master_waitrequest,           //                outgoing_master.waitrequest
		input  wire [31:0] outgoing_master_readdata,              //                               .readdata
		input  wire        outgoing_master_readdatavalid,         //                               .readdatavalid
		output wire [0:0]  outgoing_master_burstcount,            //                               .burstcount
		output wire [31:0] outgoing_master_writedata,             //                               .writedata
		output wire [26:0] outgoing_master_address,               //                               .address
		output wire        outgoing_master_write,                 //                               .write
		output wire        outgoing_master_read,                  //                               .read
		output wire [3:0]  outgoing_master_byteenable,            //                               .byteenable
		output wire        outgoing_master_debugaccess,           //                               .debugaccess
		input  wire        button_pio_external_connection_export, // button_pio_external_connection.export
		output wire        cpu0_jtag_debug_module_reset_reset,    //   cpu0_jtag_debug_module_reset.reset
		input  wire        reset_reset_n,                         //                          reset.reset_n
		input  wire        fprint_irq_0_irq_export,               //               fprint_irq_0_irq.export
		input  wire [7:0]  cpu_irq_0_s0_address,                  //                   cpu_irq_0_s0.address
		input  wire        cpu_irq_0_s0_write,                    //                               .write
		input  wire [31:0] cpu_irq_0_s0_writedata                 //                               .writedata
	);

	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_cpu0_jtag_debug_module_waitrequest;      // cpu0:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu0_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu0_jtag_debug_module_writedata;        // mm_interconnect_0:cpu0_jtag_debug_module_writedata -> cpu0:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu0_jtag_debug_module_address;          // mm_interconnect_0:cpu0_jtag_debug_module_address -> cpu0:jtag_debug_module_address
	wire         mm_interconnect_0_cpu0_jtag_debug_module_write;            // mm_interconnect_0:cpu0_jtag_debug_module_write -> cpu0:jtag_debug_module_write
	wire         mm_interconnect_0_cpu0_jtag_debug_module_read;             // mm_interconnect_0:cpu0_jtag_debug_module_read -> cpu0:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu0_jtag_debug_module_readdata;         // cpu0:jtag_debug_module_readdata -> mm_interconnect_0:cpu0_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu0_jtag_debug_module_debugaccess;      // mm_interconnect_0:cpu0_jtag_debug_module_debugaccess -> cpu0:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu0_jtag_debug_module_byteenable;       // mm_interconnect_0:cpu0_jtag_debug_module_byteenable -> cpu0:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_button_pio_s1_writedata;                 // mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	wire   [1:0] mm_interconnect_0_button_pio_s1_address;                   // mm_interconnect_0:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_0_button_pio_s1_chipselect;                // mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	wire         mm_interconnect_0_button_pio_s1_write;                     // mm_interconnect_0:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_0_button_pio_s1_readdata;                  // button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	wire         cpu0_data_master_waitrequest;                              // mm_interconnect_0:cpu0_data_master_waitrequest -> cpu0:d_waitrequest
	wire  [31:0] cpu0_data_master_writedata;                                // cpu0:d_writedata -> mm_interconnect_0:cpu0_data_master_writedata
	wire  [27:0] cpu0_data_master_address;                                  // cpu0:d_address -> mm_interconnect_0:cpu0_data_master_address
	wire         cpu0_data_master_write;                                    // cpu0:d_write -> mm_interconnect_0:cpu0_data_master_write
	wire         cpu0_data_master_read;                                     // cpu0:d_read -> mm_interconnect_0:cpu0_data_master_read
	wire  [31:0] cpu0_data_master_readdata;                                 // mm_interconnect_0:cpu0_data_master_readdata -> cpu0:d_readdata
	wire         cpu0_data_master_debugaccess;                              // cpu0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu0_data_master_debugaccess
	wire   [3:0] cpu0_data_master_byteenable;                               // cpu0:d_byteenable -> mm_interconnect_0:cpu0_data_master_byteenable
	wire  [15:0] mm_interconnect_0_timestamp_s1_writedata;                  // mm_interconnect_0:timestamp_s1_writedata -> timestamp:writedata
	wire   [3:0] mm_interconnect_0_timestamp_s1_address;                    // mm_interconnect_0:timestamp_s1_address -> timestamp:address
	wire         mm_interconnect_0_timestamp_s1_chipselect;                 // mm_interconnect_0:timestamp_s1_chipselect -> timestamp:chipselect
	wire         mm_interconnect_0_timestamp_s1_write;                      // mm_interconnect_0:timestamp_s1_write -> timestamp:write_n
	wire  [15:0] mm_interconnect_0_timestamp_s1_readdata;                   // timestamp:readdata -> mm_interconnect_0:timestamp_s1_readdata
	wire         mm_interconnect_0_out_system_bridge_s0_waitrequest;        // out_system_bridge:s0_waitrequest -> mm_interconnect_0:out_system_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_out_system_bridge_s0_burstcount;         // mm_interconnect_0:out_system_bridge_s0_burstcount -> out_system_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_writedata;          // mm_interconnect_0:out_system_bridge_s0_writedata -> out_system_bridge:s0_writedata
	wire  [26:0] mm_interconnect_0_out_system_bridge_s0_address;            // mm_interconnect_0:out_system_bridge_s0_address -> out_system_bridge:s0_address
	wire         mm_interconnect_0_out_system_bridge_s0_write;              // mm_interconnect_0:out_system_bridge_s0_write -> out_system_bridge:s0_write
	wire         mm_interconnect_0_out_system_bridge_s0_read;               // mm_interconnect_0:out_system_bridge_s0_read -> out_system_bridge:s0_read
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_readdata;           // out_system_bridge:s0_readdata -> mm_interconnect_0:out_system_bridge_s0_readdata
	wire         mm_interconnect_0_out_system_bridge_s0_debugaccess;        // mm_interconnect_0:out_system_bridge_s0_debugaccess -> out_system_bridge:s0_debugaccess
	wire         mm_interconnect_0_out_system_bridge_s0_readdatavalid;      // out_system_bridge:s0_readdatavalid -> mm_interconnect_0:out_system_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_out_system_bridge_s0_byteenable;         // mm_interconnect_0:out_system_bridge_s0_byteenable -> out_system_bridge:s0_byteenable
	wire         cpu0_instruction_master_waitrequest;                       // mm_interconnect_0:cpu0_instruction_master_waitrequest -> cpu0:i_waitrequest
	wire  [27:0] cpu0_instruction_master_address;                           // cpu0:i_address -> mm_interconnect_0:cpu0_instruction_master_address
	wire         cpu0_instruction_master_read;                              // cpu0:i_read -> mm_interconnect_0:cpu0_instruction_master_read
	wire  [31:0] cpu0_instruction_master_readdata;                          // mm_interconnect_0:cpu0_instruction_master_readdata -> cpu0:i_readdata
	wire         cpu0_instruction_master_readdatavalid;                     // mm_interconnect_0:cpu0_instruction_master_readdatavalid -> cpu0:i_readdatavalid
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire         irq_mapper_receiver0_irq;                                  // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // button_pio:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // fprint_irq_0:irq_out -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                  // cpu_irq_0:ins_irq0_irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu0_d_irq_irq;                                            // irq_mapper:sender_irq -> cpu0:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [button_pio:reset_n, cpu0:reset_n, cpu_irq_0:reset, fprint_irq_0:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpu0_reset_n_reset_bridge_in_reset_reset, out_system_bridge:reset, rst_translator:in_reset, timer:reset_n, timestamp:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [cpu0:reset_req, rst_translator:reset_req_in]

	nios_fprint_processorMonitor_cpu0 cpu0 (
		.clk                                   (philosopher_clk_in_clk),                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (cpu0_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu0_data_master_read),                                //                          .read
		.d_readdata                            (cpu0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu0_data_master_write),                               //                          .write
		.d_writedata                           (cpu0_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu0_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                      // custom_instruction_master.readra
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (27),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) out_system_bridge (
		.clk              (philosopher_clk_in_clk),                               //   clk.clk
		.reset            (rst_controller_reset_out_reset),                       // reset.reset
		.s0_waitrequest   (mm_interconnect_0_out_system_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_out_system_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_out_system_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_out_system_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_out_system_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_out_system_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_out_system_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_out_system_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_out_system_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_out_system_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (outgoing_master_waitrequest),                          //    m0.waitrequest
		.m0_readdata      (outgoing_master_readdata),                             //      .readdata
		.m0_readdatavalid (outgoing_master_readdatavalid),                        //      .readdatavalid
		.m0_burstcount    (outgoing_master_burstcount),                           //      .burstcount
		.m0_writedata     (outgoing_master_writedata),                            //      .writedata
		.m0_address       (outgoing_master_address),                              //      .address
		.m0_write         (outgoing_master_write),                                //      .write
		.m0_read          (outgoing_master_read),                                 //      .read
		.m0_byteenable    (outgoing_master_byteenable),                           //      .byteenable
		.m0_debugaccess   (outgoing_master_debugaccess)                           //      .debugaccess
	);

	nios_fprint_processorMonitor_timer timer (
		.clk        (philosopher_clk_in_clk),                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	nios_fprint_processorMonitor_jtag_uart jtag_uart (
		.clk            (philosopher_clk_in_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	nios_fprint_processorMonitor_button_pio button_pio (
		.clk        (philosopher_clk_in_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                    //                 irq.irq
	);

	fprint_irq fprint_irq_0 (
		.irq_out (irq_mapper_receiver3_irq),       // interrupt_sender.irq
		.irq     (fprint_irq_0_irq_export),        //              irq.export
		.clk     (philosopher_clk_in_clk),         //            clock.clk
		.reset   (rst_controller_reset_out_reset)  //            reset.reset
	);

	cpu_irq cpu_irq_0 (
		.avs_s0_address   (cpu_irq_0_s0_address),           //    s0.address
		.avs_s0_write     (cpu_irq_0_s0_write),             //      .write
		.avs_s0_writedata (cpu_irq_0_s0_writedata),         //      .writedata
		.clk              (philosopher_clk_in_clk),         // clock.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.ins_irq0_irq     (irq_mapper_receiver4_irq)        //  irq0.irq
	);

	nios_fprint_processorMonitor_timestamp timestamp (
		.clk        (philosopher_clk_in_clk),                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_timestamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timestamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timestamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timestamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timestamp_s1_write),     //      .write_n
		.irq        ()                                           //   irq.irq
	);

	nios_fprint_processorMonitor_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                              (philosopher_clk_in_clk),                                    //                            clk_clk.clk
		.cpu0_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpu0_reset_n_reset_bridge_in_reset.reset
		.cpu0_data_master_address                 (cpu0_data_master_address),                                  //                   cpu0_data_master.address
		.cpu0_data_master_waitrequest             (cpu0_data_master_waitrequest),                              //                                   .waitrequest
		.cpu0_data_master_byteenable              (cpu0_data_master_byteenable),                               //                                   .byteenable
		.cpu0_data_master_read                    (cpu0_data_master_read),                                     //                                   .read
		.cpu0_data_master_readdata                (cpu0_data_master_readdata),                                 //                                   .readdata
		.cpu0_data_master_write                   (cpu0_data_master_write),                                    //                                   .write
		.cpu0_data_master_writedata               (cpu0_data_master_writedata),                                //                                   .writedata
		.cpu0_data_master_debugaccess             (cpu0_data_master_debugaccess),                              //                                   .debugaccess
		.cpu0_instruction_master_address          (cpu0_instruction_master_address),                           //            cpu0_instruction_master.address
		.cpu0_instruction_master_waitrequest      (cpu0_instruction_master_waitrequest),                       //                                   .waitrequest
		.cpu0_instruction_master_read             (cpu0_instruction_master_read),                              //                                   .read
		.cpu0_instruction_master_readdata         (cpu0_instruction_master_readdata),                          //                                   .readdata
		.cpu0_instruction_master_readdatavalid    (cpu0_instruction_master_readdatavalid),                     //                                   .readdatavalid
		.button_pio_s1_address                    (mm_interconnect_0_button_pio_s1_address),                   //                      button_pio_s1.address
		.button_pio_s1_write                      (mm_interconnect_0_button_pio_s1_write),                     //                                   .write
		.button_pio_s1_readdata                   (mm_interconnect_0_button_pio_s1_readdata),                  //                                   .readdata
		.button_pio_s1_writedata                  (mm_interconnect_0_button_pio_s1_writedata),                 //                                   .writedata
		.button_pio_s1_chipselect                 (mm_interconnect_0_button_pio_s1_chipselect),                //                                   .chipselect
		.cpu0_jtag_debug_module_address           (mm_interconnect_0_cpu0_jtag_debug_module_address),          //             cpu0_jtag_debug_module.address
		.cpu0_jtag_debug_module_write             (mm_interconnect_0_cpu0_jtag_debug_module_write),            //                                   .write
		.cpu0_jtag_debug_module_read              (mm_interconnect_0_cpu0_jtag_debug_module_read),             //                                   .read
		.cpu0_jtag_debug_module_readdata          (mm_interconnect_0_cpu0_jtag_debug_module_readdata),         //                                   .readdata
		.cpu0_jtag_debug_module_writedata         (mm_interconnect_0_cpu0_jtag_debug_module_writedata),        //                                   .writedata
		.cpu0_jtag_debug_module_byteenable        (mm_interconnect_0_cpu0_jtag_debug_module_byteenable),       //                                   .byteenable
		.cpu0_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu0_jtag_debug_module_waitrequest),      //                                   .waitrequest
		.cpu0_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu0_jtag_debug_module_debugaccess),      //                                   .debugaccess
		.jtag_uart_avalon_jtag_slave_address      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                   .write
		.jtag_uart_avalon_jtag_slave_read         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                   .read
		.jtag_uart_avalon_jtag_slave_readdata     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.out_system_bridge_s0_address             (mm_interconnect_0_out_system_bridge_s0_address),            //               out_system_bridge_s0.address
		.out_system_bridge_s0_write               (mm_interconnect_0_out_system_bridge_s0_write),              //                                   .write
		.out_system_bridge_s0_read                (mm_interconnect_0_out_system_bridge_s0_read),               //                                   .read
		.out_system_bridge_s0_readdata            (mm_interconnect_0_out_system_bridge_s0_readdata),           //                                   .readdata
		.out_system_bridge_s0_writedata           (mm_interconnect_0_out_system_bridge_s0_writedata),          //                                   .writedata
		.out_system_bridge_s0_burstcount          (mm_interconnect_0_out_system_bridge_s0_burstcount),         //                                   .burstcount
		.out_system_bridge_s0_byteenable          (mm_interconnect_0_out_system_bridge_s0_byteenable),         //                                   .byteenable
		.out_system_bridge_s0_readdatavalid       (mm_interconnect_0_out_system_bridge_s0_readdatavalid),      //                                   .readdatavalid
		.out_system_bridge_s0_waitrequest         (mm_interconnect_0_out_system_bridge_s0_waitrequest),        //                                   .waitrequest
		.out_system_bridge_s0_debugaccess         (mm_interconnect_0_out_system_bridge_s0_debugaccess),        //                                   .debugaccess
		.timer_s1_address                         (mm_interconnect_0_timer_s1_address),                        //                           timer_s1.address
		.timer_s1_write                           (mm_interconnect_0_timer_s1_write),                          //                                   .write
		.timer_s1_readdata                        (mm_interconnect_0_timer_s1_readdata),                       //                                   .readdata
		.timer_s1_writedata                       (mm_interconnect_0_timer_s1_writedata),                      //                                   .writedata
		.timer_s1_chipselect                      (mm_interconnect_0_timer_s1_chipselect),                     //                                   .chipselect
		.timestamp_s1_address                     (mm_interconnect_0_timestamp_s1_address),                    //                       timestamp_s1.address
		.timestamp_s1_write                       (mm_interconnect_0_timestamp_s1_write),                      //                                   .write
		.timestamp_s1_readdata                    (mm_interconnect_0_timestamp_s1_readdata),                   //                                   .readdata
		.timestamp_s1_writedata                   (mm_interconnect_0_timestamp_s1_writedata),                  //                                   .writedata
		.timestamp_s1_chipselect                  (mm_interconnect_0_timestamp_s1_chipselect)                  //                                   .chipselect
	);

	nios_fprint_processorMonitor_irq_mapper irq_mapper (
		.clk           (philosopher_clk_in_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (cpu0_d_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (philosopher_clk_in_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
