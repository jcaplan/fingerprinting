// nios_fprint_processor1_0.v

// Generated using ACDS version 13.1 162 at 2015.06.23.14:23:19

`timescale 1 ps / 1 ps
module nios_fprint_processor1_0 (
		input  wire        philosopher_clk_in_clk,                  //             philosopher_clk_in.clk
		input  wire        outgoing_master_waitrequest,             //                outgoing_master.waitrequest
		input  wire [31:0] outgoing_master_readdata,                //                               .readdata
		input  wire        outgoing_master_readdatavalid,           //                               .readdatavalid
		output wire [0:0]  outgoing_master_burstcount,              //                               .burstcount
		output wire [31:0] outgoing_master_writedata,               //                               .writedata
		output wire [25:0] outgoing_master_address,                 //                               .address
		output wire        outgoing_master_write,                   //                               .write
		output wire        outgoing_master_read,                    //                               .read
		output wire [3:0]  outgoing_master_byteenable,              //                               .byteenable
		output wire        outgoing_master_debugaccess,             //                               .debugaccess
		input  wire        button_pio_external_connection_export,   // button_pio_external_connection.export
		input  wire        reset_reset_n,                           //                          reset.reset_n
		output wire        cpu1_jtag_debug_module_reset_reset,      //   cpu1_jtag_debug_module_reset.reset
		input  wire [7:0]  cpu1_irq_0_s0_address,                   //                  cpu1_irq_0_s0.address
		input  wire        cpu1_irq_0_s0_write,                     //                               .write
		input  wire [31:0] cpu1_irq_0_s0_writedata,                 //                               .writedata
		output wire        dma_0_irq_irq,                           //                      dma_0_irq.irq
		output wire [26:0] fingerprint_0_avalon_master_address,     //    fingerprint_0_avalon_master.address
		input  wire        fingerprint_0_avalon_master_waitrequest, //                               .waitrequest
		input  wire [31:0] fingerprint_0_avalon_master_readdata,    //                               .readdata
		output wire        fingerprint_0_avalon_master_write,       //                               .write
		output wire [31:0] fingerprint_0_avalon_master_writedata,   //                               .writedata
		output wire        fingerprint_0_avalon_master_read,        //                               .read
		input  wire [2:0]  dma_0_control_port_slave_address,        //       dma_0_control_port_slave.address
		input  wire        dma_0_control_port_slave_chipselect,     //                               .chipselect
		output wire [26:0] dma_0_control_port_slave_readdata,       //                               .readdata
		input  wire        dma_0_control_port_slave_write_n,        //                               .write_n
		input  wire [26:0] dma_0_control_port_slave_writedata,      //                               .writedata
		input  wire [7:0]  sw_reset_0_s0_address,                   //                  sw_reset_0_s0.address
		input  wire        sw_reset_0_s0_read,                      //                               .read
		output wire [31:0] sw_reset_0_s0_readdata,                  //                               .readdata
		input  wire        sw_reset_0_s0_write,                     //                               .write
		input  wire [31:0] sw_reset_0_s0_writedata,                 //                               .writedata
		output wire        sw_reset_0_s0_waitrequest,               //                               .waitrequest
		output wire        sw_reset_0_reset_source_reset            //        sw_reset_0_reset_source.reset
	);

	wire         utlb_0_fprint_waitrequest;                                                  // utlb_0:fprint_waitrequest -> Fingerprint_0:waitrequest
	wire  [31:0] utlb_0_fprint_writedata;                                                    // utlb_0:fprint_writedata -> Fingerprint_0:writedata
	wire  [26:0] utlb_0_fprint_data_address;                                                 // utlb_0:fprint_data_address -> Fingerprint_0:data_address
	wire         utlb_0_fprint_write;                                                        // utlb_0:fprint_write -> Fingerprint_0:write
	wire  [31:0] cpu1_custom_instruction_master_result;                                      // cpu1_custom_instruction_master_translator:ci_slave_result -> cpu1:E_ci_combo_result
	wire   [7:0] cpu1_custom_instruction_master_multi_n;                                     // cpu1:A_ci_multi_n -> cpu1_custom_instruction_master_translator:ci_slave_multi_n
	wire         cpu1_custom_instruction_master_writerc;                                     // cpu1:E_ci_combo_writerc -> cpu1_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] cpu1_custom_instruction_master_multi_result;                                // cpu1_custom_instruction_master_translator:ci_slave_multi_result -> cpu1:A_ci_multi_result
	wire  [31:0] cpu1_custom_instruction_master_multi_dataa;                                 // cpu1:A_ci_multi_dataa -> cpu1_custom_instruction_master_translator:ci_slave_multi_dataa
	wire  [31:0] cpu1_custom_instruction_master_dataa;                                       // cpu1:E_ci_combo_dataa -> cpu1_custom_instruction_master_translator:ci_slave_dataa
	wire  [31:0] cpu1_custom_instruction_master_multi_datab;                                 // cpu1:A_ci_multi_datab -> cpu1_custom_instruction_master_translator:ci_slave_multi_datab
	wire         cpu1_custom_instruction_master_readra;                                      // cpu1:E_ci_combo_readra -> cpu1_custom_instruction_master_translator:ci_slave_readra
	wire         cpu1_custom_instruction_master_reset;                                       // cpu1:A_ci_multi_reset -> cpu1_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] cpu1_custom_instruction_master_datab;                                       // cpu1:E_ci_combo_datab -> cpu1_custom_instruction_master_translator:ci_slave_datab
	wire         cpu1_custom_instruction_master_readrb;                                      // cpu1:E_ci_combo_readrb -> cpu1_custom_instruction_master_translator:ci_slave_readrb
	wire         cpu1_custom_instruction_master_multi_readra;                                // cpu1:A_ci_multi_readra -> cpu1_custom_instruction_master_translator:ci_slave_multi_readra
	wire         cpu1_custom_instruction_master_multi_readrb;                                // cpu1:A_ci_multi_readrb -> cpu1_custom_instruction_master_translator:ci_slave_multi_readrb
	wire   [4:0] cpu1_custom_instruction_master_b;                                           // cpu1:E_ci_combo_b -> cpu1_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] cpu1_custom_instruction_master_c;                                           // cpu1:E_ci_combo_c -> cpu1_custom_instruction_master_translator:ci_slave_c
	wire         cpu1_custom_instruction_master_clk_en;                                      // cpu1:A_ci_multi_clk_en -> cpu1_custom_instruction_master_translator:ci_slave_multi_clken
	wire         cpu1_custom_instruction_master_done;                                        // cpu1_custom_instruction_master_translator:ci_slave_multi_done -> cpu1:A_ci_multi_done
	wire   [4:0] cpu1_custom_instruction_master_a;                                           // cpu1:E_ci_combo_a -> cpu1_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] cpu1_custom_instruction_master_n;                                           // cpu1:E_ci_combo_n -> cpu1_custom_instruction_master_translator:ci_slave_n
	wire         cpu1_custom_instruction_master_multi_writerc;                               // cpu1:A_ci_multi_writerc -> cpu1_custom_instruction_master_translator:ci_slave_multi_writerc
	wire         cpu1_custom_instruction_master_clk;                                         // cpu1:A_ci_multi_clock -> cpu1_custom_instruction_master_translator:ci_slave_multi_clk
	wire         cpu1_custom_instruction_master_reset_req;                                   // cpu1:A_ci_multi_reset_req -> cpu1_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] cpu1_custom_instruction_master_multi_c;                                     // cpu1:A_ci_multi_c -> cpu1_custom_instruction_master_translator:ci_slave_multi_c
	wire   [4:0] cpu1_custom_instruction_master_multi_b;                                     // cpu1:A_ci_multi_b -> cpu1_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] cpu1_custom_instruction_master_multi_a;                                     // cpu1:A_ci_multi_a -> cpu1_custom_instruction_master_translator:ci_slave_multi_a
	wire         cpu1_custom_instruction_master_start;                                       // cpu1:A_ci_multi_start -> cpu1_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] cpu1_custom_instruction_master_translator_comb_ci_master_result;            // cpu1_custom_instruction_master_comb_xconnect:ci_slave_result -> cpu1_custom_instruction_master_translator:comb_ci_master_result
	wire   [4:0] cpu1_custom_instruction_master_translator_comb_ci_master_b;                 // cpu1_custom_instruction_master_translator:comb_ci_master_b -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_b
	wire   [4:0] cpu1_custom_instruction_master_translator_comb_ci_master_c;                 // cpu1_custom_instruction_master_translator:comb_ci_master_c -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_c
	wire  [31:0] cpu1_custom_instruction_master_translator_comb_ci_master_dataa;             // cpu1_custom_instruction_master_translator:comb_ci_master_dataa -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire   [4:0] cpu1_custom_instruction_master_translator_comb_ci_master_a;                 // cpu1_custom_instruction_master_translator:comb_ci_master_a -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_a
	wire         cpu1_custom_instruction_master_translator_comb_ci_master_readra;            // cpu1_custom_instruction_master_translator:comb_ci_master_readra -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [7:0] cpu1_custom_instruction_master_translator_comb_ci_master_n;                 // cpu1_custom_instruction_master_translator:comb_ci_master_n -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_n
	wire         cpu1_custom_instruction_master_translator_comb_ci_master_writerc;           // cpu1_custom_instruction_master_translator:comb_ci_master_writerc -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire  [31:0] cpu1_custom_instruction_master_translator_comb_ci_master_datab;             // cpu1_custom_instruction_master_translator:comb_ci_master_datab -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] cpu1_custom_instruction_master_translator_comb_ci_master_ipending;          // cpu1_custom_instruction_master_translator:comb_ci_master_ipending -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire         cpu1_custom_instruction_master_translator_comb_ci_master_readrb;            // cpu1_custom_instruction_master_translator:comb_ci_master_readrb -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire         cpu1_custom_instruction_master_translator_comb_ci_master_estatus;           // cpu1_custom_instruction_master_translator:comb_ci_master_estatus -> cpu1_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] cpu1_custom_instruction_master_comb_xconnect_ci_master0_result;             // cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpu1_custom_instruction_master_comb_xconnect:ci_master0_result
	wire   [4:0] cpu1_custom_instruction_master_comb_xconnect_ci_master0_b;                  // cpu1_custom_instruction_master_comb_xconnect:ci_master0_b -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire   [4:0] cpu1_custom_instruction_master_comb_xconnect_ci_master0_c;                  // cpu1_custom_instruction_master_comb_xconnect:ci_master0_c -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire  [31:0] cpu1_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // cpu1_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire   [4:0] cpu1_custom_instruction_master_comb_xconnect_ci_master0_a;                  // cpu1_custom_instruction_master_comb_xconnect:ci_master0_a -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire         cpu1_custom_instruction_master_comb_xconnect_ci_master0_readra;             // cpu1_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [7:0] cpu1_custom_instruction_master_comb_xconnect_ci_master0_n;                  // cpu1_custom_instruction_master_comb_xconnect:ci_master0_n -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire         cpu1_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // cpu1_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire  [31:0] cpu1_custom_instruction_master_comb_xconnect_ci_master0_datab;              // cpu1_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] cpu1_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // cpu1_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire         cpu1_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // cpu1_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire         cpu1_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // cpu1_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpu1_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu1_custom_instruction_master_comb_slave_translator0_ci_master_result;     // nios_custom_instr_floating_point_2_0:s1_result -> cpu1_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] cpu1_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // cpu1_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s1_dataa
	wire   [3:0] cpu1_custom_instruction_master_comb_slave_translator0_ci_master_n;          // cpu1_custom_instruction_master_comb_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s1_n
	wire  [31:0] cpu1_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // cpu1_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s1_datab
	wire  [31:0] cpu1_custom_instruction_master_translator_multi_ci_master_result;           // cpu1_custom_instruction_master_multi_xconnect:ci_slave_result -> cpu1_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] cpu1_custom_instruction_master_translator_multi_ci_master_b;                // cpu1_custom_instruction_master_translator:multi_ci_master_b -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] cpu1_custom_instruction_master_translator_multi_ci_master_c;                // cpu1_custom_instruction_master_translator:multi_ci_master_c -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] cpu1_custom_instruction_master_translator_multi_ci_master_a;                // cpu1_custom_instruction_master_translator:multi_ci_master_a -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_clk_en;           // cpu1_custom_instruction_master_translator:multi_ci_master_clken -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_done;             // cpu1_custom_instruction_master_multi_xconnect:ci_slave_done -> cpu1_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] cpu1_custom_instruction_master_translator_multi_ci_master_n;                // cpu1_custom_instruction_master_translator:multi_ci_master_n -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_writerc;          // cpu1_custom_instruction_master_translator:multi_ci_master_writerc -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_clk;              // cpu1_custom_instruction_master_translator:multi_ci_master_clk -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_reset_req;        // cpu1_custom_instruction_master_translator:multi_ci_master_reset_req -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_start;            // cpu1_custom_instruction_master_translator:multi_ci_master_start -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] cpu1_custom_instruction_master_translator_multi_ci_master_dataa;            // cpu1_custom_instruction_master_translator:multi_ci_master_dataa -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_readra;           // cpu1_custom_instruction_master_translator:multi_ci_master_readra -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_reset;            // cpu1_custom_instruction_master_translator:multi_ci_master_reset -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] cpu1_custom_instruction_master_translator_multi_ci_master_datab;            // cpu1_custom_instruction_master_translator:multi_ci_master_datab -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         cpu1_custom_instruction_master_translator_multi_ci_master_readrb;           // cpu1_custom_instruction_master_translator:multi_ci_master_readrb -> cpu1_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] cpu1_custom_instruction_master_multi_xconnect_ci_master0_result;            // cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpu1_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] cpu1_custom_instruction_master_multi_xconnect_ci_master0_b;                 // cpu1_custom_instruction_master_multi_xconnect:ci_master0_b -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] cpu1_custom_instruction_master_multi_xconnect_ci_master0_c;                 // cpu1_custom_instruction_master_multi_xconnect:ci_master0_c -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_done;              // cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpu1_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // cpu1_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] cpu1_custom_instruction_master_multi_xconnect_ci_master0_a;                 // cpu1_custom_instruction_master_multi_xconnect:ci_master0_a -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] cpu1_custom_instruction_master_multi_xconnect_ci_master0_n;                 // cpu1_custom_instruction_master_multi_xconnect:ci_master0_n -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // cpu1_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] cpu1_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // cpu1_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_clk;               // cpu1_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // cpu1_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_start;             // cpu1_custom_instruction_master_multi_xconnect:ci_master0_start -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] cpu1_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // cpu1_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_readra;            // cpu1_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_reset;             // cpu1_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] cpu1_custom_instruction_master_multi_xconnect_ci_master0_datab;             // cpu1_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // cpu1_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         cpu1_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // cpu1_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpu1_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] cpu1_custom_instruction_master_multi_slave_translator0_ci_master_result;    // nios_custom_instr_floating_point_2_0:s2_result -> cpu1_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         cpu1_custom_instruction_master_multi_slave_translator0_ci_master_start;     // cpu1_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_2_0:s2_start
	wire  [31:0] cpu1_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // cpu1_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s2_dataa
	wire         cpu1_custom_instruction_master_multi_slave_translator0_ci_master_done;      // nios_custom_instr_floating_point_2_0:s2_done -> cpu1_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         cpu1_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // cpu1_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_2_0:s2_clk_en
	wire   [2:0] cpu1_custom_instruction_master_multi_slave_translator0_ci_master_n;         // cpu1_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s2_n
	wire         cpu1_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // cpu1_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_2_0:s2_reset
	wire  [31:0] cpu1_custom_instruction_master_multi_slave_translator0_ci_master_datab;     // cpu1_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s2_datab
	wire         cpu1_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // cpu1_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_2_0:s2_clk
	wire         cpu1_custom_instruction_master_multi_slave_translator0_ci_master_reset_req; // cpu1_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> nios_custom_instr_floating_point_2_0:s2_reset_req
	wire         dma_0_read_master_waitrequest;                                              // mm_interconnect_0:dma_0_read_master_waitrequest -> dma_0:read_waitrequest
	wire  [26:0] dma_0_read_master_address;                                                  // dma_0:read_address -> mm_interconnect_0:dma_0_read_master_address
	wire         dma_0_read_master_chipselect;                                               // dma_0:read_chipselect -> mm_interconnect_0:dma_0_read_master_chipselect
	wire         dma_0_read_master_read;                                                     // dma_0:read_read_n -> mm_interconnect_0:dma_0_read_master_read
	wire  [31:0] dma_0_read_master_readdata;                                                 // mm_interconnect_0:dma_0_read_master_readdata -> dma_0:read_readdata
	wire         dma_0_read_master_readdatavalid;                                            // mm_interconnect_0:dma_0_read_master_readdatavalid -> dma_0:read_readdatavalid
	wire  [31:0] mm_interconnect_0_scratchpad_1_s1_writedata;                                // mm_interconnect_0:scratchpad_1_s1_writedata -> scratchpad_1:writedata
	wire  [11:0] mm_interconnect_0_scratchpad_1_s1_address;                                  // mm_interconnect_0:scratchpad_1_s1_address -> scratchpad_1:address
	wire         mm_interconnect_0_scratchpad_1_s1_chipselect;                               // mm_interconnect_0:scratchpad_1_s1_chipselect -> scratchpad_1:chipselect
	wire         mm_interconnect_0_scratchpad_1_s1_clken;                                    // mm_interconnect_0:scratchpad_1_s1_clken -> scratchpad_1:clken
	wire         mm_interconnect_0_scratchpad_1_s1_write;                                    // mm_interconnect_0:scratchpad_1_s1_write -> scratchpad_1:write
	wire  [31:0] mm_interconnect_0_scratchpad_1_s1_readdata;                                 // scratchpad_1:readdata -> mm_interconnect_0:scratchpad_1_s1_readdata
	wire   [3:0] mm_interconnect_0_scratchpad_1_s1_byteenable;                               // mm_interconnect_0:scratchpad_1_s1_byteenable -> scratchpad_1:byteenable
	wire         dma_0_write_master_waitrequest;                                             // mm_interconnect_0:dma_0_write_master_waitrequest -> dma_0:write_waitrequest
	wire  [31:0] dma_0_write_master_writedata;                                               // dma_0:write_writedata -> mm_interconnect_0:dma_0_write_master_writedata
	wire  [26:0] dma_0_write_master_address;                                                 // dma_0:write_address -> mm_interconnect_0:dma_0_write_master_address
	wire         dma_0_write_master_chipselect;                                              // dma_0:write_chipselect -> mm_interconnect_0:dma_0_write_master_chipselect
	wire         dma_0_write_master_write;                                                   // dma_0:write_write_n -> mm_interconnect_0:dma_0_write_master_write
	wire   [3:0] dma_0_write_master_byteenable;                                              // dma_0:write_byteenable -> mm_interconnect_0:dma_0_write_master_byteenable
	wire         mm_interconnect_0_out_system_bridge_s0_waitrequest;                         // out_system_bridge:s0_waitrequest -> mm_interconnect_0:out_system_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_out_system_bridge_s0_burstcount;                          // mm_interconnect_0:out_system_bridge_s0_burstcount -> out_system_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_writedata;                           // mm_interconnect_0:out_system_bridge_s0_writedata -> out_system_bridge:s0_writedata
	wire  [25:0] mm_interconnect_0_out_system_bridge_s0_address;                             // mm_interconnect_0:out_system_bridge_s0_address -> out_system_bridge:s0_address
	wire         mm_interconnect_0_out_system_bridge_s0_write;                               // mm_interconnect_0:out_system_bridge_s0_write -> out_system_bridge:s0_write
	wire         mm_interconnect_0_out_system_bridge_s0_read;                                // mm_interconnect_0:out_system_bridge_s0_read -> out_system_bridge:s0_read
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_readdata;                            // out_system_bridge:s0_readdata -> mm_interconnect_0:out_system_bridge_s0_readdata
	wire         mm_interconnect_0_out_system_bridge_s0_debugaccess;                         // mm_interconnect_0:out_system_bridge_s0_debugaccess -> out_system_bridge:s0_debugaccess
	wire         mm_interconnect_0_out_system_bridge_s0_readdatavalid;                       // out_system_bridge:s0_readdatavalid -> mm_interconnect_0:out_system_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_out_system_bridge_s0_byteenable;                          // mm_interconnect_0:out_system_bridge_s0_byteenable -> out_system_bridge:s0_byteenable
	wire  [31:0] mm_interconnect_0_scratchpad_0_s1_writedata;                                // mm_interconnect_0:scratchpad_0_s1_writedata -> scratchpad_0:writedata
	wire  [11:0] mm_interconnect_0_scratchpad_0_s1_address;                                  // mm_interconnect_0:scratchpad_0_s1_address -> scratchpad_0:address
	wire         mm_interconnect_0_scratchpad_0_s1_chipselect;                               // mm_interconnect_0:scratchpad_0_s1_chipselect -> scratchpad_0:chipselect
	wire         mm_interconnect_0_scratchpad_0_s1_clken;                                    // mm_interconnect_0:scratchpad_0_s1_clken -> scratchpad_0:clken
	wire         mm_interconnect_0_scratchpad_0_s1_write;                                    // mm_interconnect_0:scratchpad_0_s1_write -> scratchpad_0:write
	wire  [31:0] mm_interconnect_0_scratchpad_0_s1_readdata;                                 // scratchpad_0:readdata -> mm_interconnect_0:scratchpad_0_s1_readdata
	wire   [3:0] mm_interconnect_0_scratchpad_0_s1_byteenable;                               // mm_interconnect_0:scratchpad_0_s1_byteenable -> scratchpad_0:byteenable
	wire         utlb_0_avalon_master_waitrequest;                                           // mm_interconnect_0:utlb_0_avalon_master_waitrequest -> utlb_0:avm_waitrequest
	wire  [26:0] utlb_0_avalon_master_address;                                               // utlb_0:avm_address -> mm_interconnect_0:utlb_0_avalon_master_address
	wire  [31:0] utlb_0_avalon_master_writedata;                                             // utlb_0:avm_writedata -> mm_interconnect_0:utlb_0_avalon_master_writedata
	wire         utlb_0_avalon_master_write;                                                 // utlb_0:avm_write -> mm_interconnect_0:utlb_0_avalon_master_write
	wire         utlb_0_avalon_master_read;                                                  // utlb_0:avm_read -> mm_interconnect_0:utlb_0_avalon_master_read
	wire  [31:0] utlb_0_avalon_master_readdata;                                              // mm_interconnect_0:utlb_0_avalon_master_readdata -> utlb_0:avm_readdata
	wire   [3:0] utlb_0_avalon_master_byteenable;                                            // utlb_0:avm_byteenable -> mm_interconnect_0:utlb_0_avalon_master_byteenable
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;                  // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;                    // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;                      // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;                   // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;                        // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                         // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;                     // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_utlb_0_avalon_slave_waitrequest;                          // utlb_0:avs_waitrequest -> mm_interconnect_1:utlb_0_avalon_slave_waitrequest
	wire  [31:0] mm_interconnect_1_utlb_0_avalon_slave_writedata;                            // mm_interconnect_1:utlb_0_avalon_slave_writedata -> utlb_0:avs_writedata
	wire  [26:0] mm_interconnect_1_utlb_0_avalon_slave_address;                              // mm_interconnect_1:utlb_0_avalon_slave_address -> utlb_0:avs_address
	wire         mm_interconnect_1_utlb_0_avalon_slave_write;                                // mm_interconnect_1:utlb_0_avalon_slave_write -> utlb_0:avs_write
	wire         mm_interconnect_1_utlb_0_avalon_slave_read;                                 // mm_interconnect_1:utlb_0_avalon_slave_read -> utlb_0:avs_read
	wire  [31:0] mm_interconnect_1_utlb_0_avalon_slave_readdata;                             // utlb_0:avs_readdata -> mm_interconnect_1:utlb_0_avalon_slave_readdata
	wire   [3:0] mm_interconnect_1_utlb_0_avalon_slave_byteenable;                           // mm_interconnect_1:utlb_0_avalon_slave_byteenable -> utlb_0:avs_byteenable
	wire         cpu1_data_master_waitrequest;                                               // mm_interconnect_1:cpu1_data_master_waitrequest -> cpu1:d_waitrequest
	wire  [31:0] cpu1_data_master_writedata;                                                 // cpu1:d_writedata -> mm_interconnect_1:cpu1_data_master_writedata
	wire  [27:0] cpu1_data_master_address;                                                   // cpu1:d_address -> mm_interconnect_1:cpu1_data_master_address
	wire         cpu1_data_master_write;                                                     // cpu1:d_write -> mm_interconnect_1:cpu1_data_master_write
	wire         cpu1_data_master_read;                                                      // cpu1:d_read -> mm_interconnect_1:cpu1_data_master_read
	wire  [31:0] cpu1_data_master_readdata;                                                  // mm_interconnect_1:cpu1_data_master_readdata -> cpu1:d_readdata
	wire         cpu1_data_master_debugaccess;                                               // cpu1:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_1:cpu1_data_master_debugaccess
	wire   [3:0] cpu1_data_master_byteenable;                                                // cpu1:d_byteenable -> mm_interconnect_1:cpu1_data_master_byteenable
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                                       // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                                         // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_chipselect;                                      // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_1_timer_s1_write;                                           // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                                        // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire         mm_interconnect_1_utlb_0_ctrl_reg_waitrequest;                              // utlb_0:avs_ctrl_reg_waitrequest -> mm_interconnect_1:utlb_0_ctrl_reg_waitrequest
	wire  [31:0] mm_interconnect_1_utlb_0_ctrl_reg_writedata;                                // mm_interconnect_1:utlb_0_ctrl_reg_writedata -> utlb_0:avs_ctrl_reg_writedata
	wire   [7:0] mm_interconnect_1_utlb_0_ctrl_reg_address;                                  // mm_interconnect_1:utlb_0_ctrl_reg_address -> utlb_0:avs_ctrl_reg_address
	wire         mm_interconnect_1_utlb_0_ctrl_reg_write;                                    // mm_interconnect_1:utlb_0_ctrl_reg_write -> utlb_0:avs_ctrl_reg_write
	wire         mm_interconnect_1_utlb_0_ctrl_reg_read;                                     // mm_interconnect_1:utlb_0_ctrl_reg_read -> utlb_0:avs_ctrl_reg_read
	wire  [31:0] mm_interconnect_1_utlb_0_ctrl_reg_readdata;                                 // utlb_0:avs_ctrl_reg_readdata -> mm_interconnect_1:utlb_0_ctrl_reg_readdata
	wire         cpu1_instruction_master_waitrequest;                                        // mm_interconnect_1:cpu1_instruction_master_waitrequest -> cpu1:i_waitrequest
	wire  [27:0] cpu1_instruction_master_address;                                            // cpu1:i_address -> mm_interconnect_1:cpu1_instruction_master_address
	wire         cpu1_instruction_master_read;                                               // cpu1:i_read -> mm_interconnect_1:cpu1_instruction_master_read
	wire  [31:0] cpu1_instruction_master_readdata;                                           // mm_interconnect_1:cpu1_instruction_master_readdata -> cpu1:i_readdata
	wire         cpu1_instruction_master_readdatavalid;                                      // mm_interconnect_1:cpu1_instruction_master_readdatavalid -> cpu1:i_readdatavalid
	wire         mm_interconnect_1_fingerprint_0_avalon_slave_0_waitrequest;                 // Fingerprint_0:slave_waitrequest -> mm_interconnect_1:Fingerprint_0_avalon_slave_0_waitrequest
	wire  [31:0] mm_interconnect_1_fingerprint_0_avalon_slave_0_writedata;                   // mm_interconnect_1:Fingerprint_0_avalon_slave_0_writedata -> Fingerprint_0:slave_spr_dat_i
	wire   [7:0] mm_interconnect_1_fingerprint_0_avalon_slave_0_address;                     // mm_interconnect_1:Fingerprint_0_avalon_slave_0_address -> Fingerprint_0:slave_spr_addr
	wire         mm_interconnect_1_fingerprint_0_avalon_slave_0_write;                       // mm_interconnect_1:Fingerprint_0_avalon_slave_0_write -> Fingerprint_0:slave_spr_write
	wire         mm_interconnect_1_fingerprint_0_avalon_slave_0_read;                        // mm_interconnect_1:Fingerprint_0_avalon_slave_0_read -> Fingerprint_0:slave_spr_read
	wire  [31:0] mm_interconnect_1_fingerprint_0_avalon_slave_0_readdata;                    // Fingerprint_0:slave_spr_dat_o -> mm_interconnect_1:Fingerprint_0_avalon_slave_0_readdata
	wire  [15:0] mm_interconnect_1_timestamp_s1_writedata;                                   // mm_interconnect_1:timestamp_s1_writedata -> timestamp:writedata
	wire   [3:0] mm_interconnect_1_timestamp_s1_address;                                     // mm_interconnect_1:timestamp_s1_address -> timestamp:address
	wire         mm_interconnect_1_timestamp_s1_chipselect;                                  // mm_interconnect_1:timestamp_s1_chipselect -> timestamp:chipselect
	wire         mm_interconnect_1_timestamp_s1_write;                                       // mm_interconnect_1:timestamp_s1_write -> timestamp:write_n
	wire  [15:0] mm_interconnect_1_timestamp_s1_readdata;                                    // timestamp:readdata -> mm_interconnect_1:timestamp_s1_readdata
	wire         mm_interconnect_1_cpu1_jtag_debug_module_waitrequest;                       // cpu1:jtag_debug_module_waitrequest -> mm_interconnect_1:cpu1_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_1_cpu1_jtag_debug_module_writedata;                         // mm_interconnect_1:cpu1_jtag_debug_module_writedata -> cpu1:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_1_cpu1_jtag_debug_module_address;                           // mm_interconnect_1:cpu1_jtag_debug_module_address -> cpu1:jtag_debug_module_address
	wire         mm_interconnect_1_cpu1_jtag_debug_module_write;                             // mm_interconnect_1:cpu1_jtag_debug_module_write -> cpu1:jtag_debug_module_write
	wire         mm_interconnect_1_cpu1_jtag_debug_module_read;                              // mm_interconnect_1:cpu1_jtag_debug_module_read -> cpu1:jtag_debug_module_read
	wire  [31:0] mm_interconnect_1_cpu1_jtag_debug_module_readdata;                          // cpu1:jtag_debug_module_readdata -> mm_interconnect_1:cpu1_jtag_debug_module_readdata
	wire         mm_interconnect_1_cpu1_jtag_debug_module_debugaccess;                       // mm_interconnect_1:cpu1_jtag_debug_module_debugaccess -> cpu1:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_1_cpu1_jtag_debug_module_byteenable;                        // mm_interconnect_1:cpu1_jtag_debug_module_byteenable -> cpu1:jtag_debug_module_byteenable
	wire         irq_mapper_receiver0_irq;                                                   // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                   // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                   // button_pio:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                   // cpu_irq_0:ins_irq0_irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu1_d_irq_irq;                                                             // irq_mapper:sender_irq -> cpu1:d_irq
	wire         rst_controller_reset_out_reset;                                             // rst_controller:reset_out -> [Fingerprint_0:rst, button_pio:reset_n, cpu1:reset_n, cpu_irq_0:reset, dma_0:system_reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:dma_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:cpu1_reset_n_reset_bridge_in_reset_reset, out_system_bridge:reset, rst_translator:in_reset, scratchpad_0:reset, scratchpad_1:reset, timer:reset_n, timestamp:reset_n, utlb_0:reset]
	wire         rst_controller_reset_out_reset_req;                                         // rst_controller:reset_req -> [cpu1:reset_req, rst_translator:reset_req_in, scratchpad_0:reset_req, scratchpad_1:reset_req]

	nios_fprint_processor1_0_cpu1 cpu1 (
		.clk                                   (philosopher_clk_in_clk),                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (cpu1_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu1_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu1_data_master_read),                                //                          .read
		.d_readdata                            (cpu1_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu1_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu1_data_master_write),                               //                          .write
		.d_writedata                           (cpu1_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu1_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu1_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu1_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu1_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu1_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu1_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu1_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu1_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_1_cpu1_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_1_cpu1_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_1_cpu1_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_1_cpu1_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_1_cpu1_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_1_cpu1_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_1_cpu1_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_1_cpu1_jtag_debug_module_writedata),   //                          .writedata
		.A_ci_multi_done                       (cpu1_custom_instruction_master_done),                  // custom_instruction_master.done
		.A_ci_multi_result                     (cpu1_custom_instruction_master_multi_result),          //                          .multi_result
		.A_ci_multi_a                          (cpu1_custom_instruction_master_multi_a),               //                          .multi_a
		.A_ci_multi_b                          (cpu1_custom_instruction_master_multi_b),               //                          .multi_b
		.A_ci_multi_c                          (cpu1_custom_instruction_master_multi_c),               //                          .multi_c
		.A_ci_multi_clk_en                     (cpu1_custom_instruction_master_clk_en),                //                          .clk_en
		.A_ci_multi_clock                      (cpu1_custom_instruction_master_clk),                   //                          .clk
		.A_ci_multi_reset                      (cpu1_custom_instruction_master_reset),                 //                          .reset
		.A_ci_multi_reset_req                  (cpu1_custom_instruction_master_reset_req),             //                          .reset_req
		.A_ci_multi_dataa                      (cpu1_custom_instruction_master_multi_dataa),           //                          .multi_dataa
		.A_ci_multi_datab                      (cpu1_custom_instruction_master_multi_datab),           //                          .multi_datab
		.A_ci_multi_n                          (cpu1_custom_instruction_master_multi_n),               //                          .multi_n
		.A_ci_multi_readra                     (cpu1_custom_instruction_master_multi_readra),          //                          .multi_readra
		.A_ci_multi_readrb                     (cpu1_custom_instruction_master_multi_readrb),          //                          .multi_readrb
		.A_ci_multi_start                      (cpu1_custom_instruction_master_start),                 //                          .start
		.A_ci_multi_writerc                    (cpu1_custom_instruction_master_multi_writerc),         //                          .multi_writerc
		.E_ci_combo_result                     (cpu1_custom_instruction_master_result),                //                          .result
		.E_ci_combo_a                          (cpu1_custom_instruction_master_a),                     //                          .a
		.E_ci_combo_b                          (cpu1_custom_instruction_master_b),                     //                          .b
		.E_ci_combo_c                          (cpu1_custom_instruction_master_c),                     //                          .c
		.E_ci_combo_dataa                      (cpu1_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_combo_datab                      (cpu1_custom_instruction_master_datab),                 //                          .datab
		.E_ci_combo_n                          (cpu1_custom_instruction_master_n),                     //                          .n
		.E_ci_combo_readra                     (cpu1_custom_instruction_master_readra),                //                          .readra
		.E_ci_combo_readrb                     (cpu1_custom_instruction_master_readrb),                //                          .readrb
		.E_ci_combo_writerc                    (cpu1_custom_instruction_master_writerc)                //                          .writerc
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (26),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) out_system_bridge (
		.clk              (philosopher_clk_in_clk),                               //   clk.clk
		.reset            (rst_controller_reset_out_reset),                       // reset.reset
		.s0_waitrequest   (mm_interconnect_0_out_system_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_out_system_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_out_system_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_out_system_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_out_system_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_out_system_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_out_system_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_out_system_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_out_system_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_out_system_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (outgoing_master_waitrequest),                          //    m0.waitrequest
		.m0_readdata      (outgoing_master_readdata),                             //      .readdata
		.m0_readdatavalid (outgoing_master_readdatavalid),                        //      .readdatavalid
		.m0_burstcount    (outgoing_master_burstcount),                           //      .burstcount
		.m0_writedata     (outgoing_master_writedata),                            //      .writedata
		.m0_address       (outgoing_master_address),                              //      .address
		.m0_write         (outgoing_master_write),                                //      .write
		.m0_read          (outgoing_master_read),                                 //      .read
		.m0_byteenable    (outgoing_master_byteenable),                           //      .byteenable
		.m0_debugaccess   (outgoing_master_debugaccess)                           //      .debugaccess
	);

	nios_fprint_processor1_0_timer timer (
		.clk        (philosopher_clk_in_clk),                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	nios_fprint_processor1_0_jtag_uart jtag_uart (
		.clk            (philosopher_clk_in_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	nios_fprint_processor1_0_button_pio button_pio (
		.clk        (philosopher_clk_in_clk),                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (),                                      //                  s1.address
		.write_n    (),                                      //                    .write_n
		.writedata  (),                                      //                    .writedata
		.chipselect (),                                      //                    .chipselect
		.readdata   (),                                      //                    .readdata
		.in_port    (button_pio_external_connection_export), // external_connection.export
		.irq        (irq_mapper_receiver2_irq)               //                 irq.irq
	);

	cpu_irq cpu_irq_0 (
		.avs_s0_address   (cpu1_irq_0_s0_address),          //    s0.address
		.avs_s0_write     (cpu1_irq_0_s0_write),            //      .write
		.avs_s0_writedata (cpu1_irq_0_s0_writedata),        //      .writedata
		.clk              (philosopher_clk_in_clk),         // clock.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.ins_irq0_irq     (irq_mapper_receiver3_irq)        //  irq0.irq
	);

	nios_fprint_processor1_0_timestamp timestamp (
		.clk        (philosopher_clk_in_clk),                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_1_timestamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timestamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timestamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timestamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timestamp_s1_write),     //      .write_n
		.irq        ()                                           //   irq.irq
	);

	crc_fingerprint #(
		.CORE_ID (1)
	) fingerprint_0 (
		.clk                (philosopher_clk_in_clk),                                     //          clock.clk
		.slave_spr_addr     (mm_interconnect_1_fingerprint_0_avalon_slave_0_address),     // avalon_slave_0.address
		.slave_spr_dat_i    (mm_interconnect_1_fingerprint_0_avalon_slave_0_writedata),   //               .writedata
		.slave_spr_dat_o    (mm_interconnect_1_fingerprint_0_avalon_slave_0_readdata),    //               .readdata
		.slave_spr_read     (mm_interconnect_1_fingerprint_0_avalon_slave_0_read),        //               .read
		.slave_spr_write    (mm_interconnect_1_fingerprint_0_avalon_slave_0_write),       //               .write
		.slave_waitrequest  (mm_interconnect_1_fingerprint_0_avalon_slave_0_waitrequest), //               .waitrequest
		.master_address     (fingerprint_0_avalon_master_address),                        //  avalon_master.address
		.master_waitrequest (fingerprint_0_avalon_master_waitrequest),                    //               .waitrequest
		.master_readdata    (fingerprint_0_avalon_master_readdata),                       //               .readdata
		.master_write       (fingerprint_0_avalon_master_write),                          //               .write
		.master_writedata   (fingerprint_0_avalon_master_writedata),                      //               .writedata
		.master_read        (fingerprint_0_avalon_master_read),                           //               .read
		.rst                (rst_controller_reset_out_reset),                             //     reset_sink.reset
		.waitrequest        (utlb_0_fprint_waitrequest),                                  // fprint_conduit.export
		.data_address       (utlb_0_fprint_data_address),                                 //               .export
		.writedata          (utlb_0_fprint_writedata),                                    //               .export
		.write              (utlb_0_fprint_write)                                         //               .export
	);

	nios_fprint_processor1_0_scratchpad_0 scratchpad_0 (
		.clk        (philosopher_clk_in_clk),                       //   clk1.clk
		.address    (mm_interconnect_0_scratchpad_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_scratchpad_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_scratchpad_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_scratchpad_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_scratchpad_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_scratchpad_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_scratchpad_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)            //       .reset_req
	);

	nios_fprint_processor1_0_dma_0 dma_0 (
		.clk                (philosopher_clk_in_clk),              //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),     //              reset.reset_n
		.dma_ctl_address    (dma_0_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (dma_0_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (dma_0_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (dma_0_control_port_slave_write_n),    //                   .write_n
		.dma_ctl_writedata  (dma_0_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (dma_0_irq_irq),                       //                irq.irq
		.read_address       (dma_0_read_master_address),           //        read_master.address
		.read_chipselect    (dma_0_read_master_chipselect),        //                   .chipselect
		.read_read_n        (dma_0_read_master_read),              //                   .read_n
		.read_readdata      (dma_0_read_master_readdata),          //                   .readdata
		.read_readdatavalid (dma_0_read_master_readdatavalid),     //                   .readdatavalid
		.read_waitrequest   (dma_0_read_master_waitrequest),       //                   .waitrequest
		.write_address      (dma_0_write_master_address),          //       write_master.address
		.write_chipselect   (dma_0_write_master_chipselect),       //                   .chipselect
		.write_waitrequest  (dma_0_write_master_waitrequest),      //                   .waitrequest
		.write_write_n      (dma_0_write_master_write),            //                   .write_n
		.write_writedata    (dma_0_write_master_writedata),        //                   .writedata
		.write_byteenable   (dma_0_write_master_byteenable)        //                   .byteenable
	);

	fulltlb #(
		.tagwidth        (15),
		.addresswidth    (27),
		.numentries      (4),
		.datawidth       (32),
		.byteenablewidth (4)
	) utlb_0 (
		.avs_ctrl_reg_address     (mm_interconnect_1_utlb_0_ctrl_reg_address),         //      ctrl_reg.address
		.avs_ctrl_reg_writedata   (mm_interconnect_1_utlb_0_ctrl_reg_writedata),       //              .writedata
		.avs_ctrl_reg_write       (mm_interconnect_1_utlb_0_ctrl_reg_write),           //              .write
		.avs_ctrl_reg_read        (mm_interconnect_1_utlb_0_ctrl_reg_read),            //              .read
		.avs_ctrl_reg_readdata    (mm_interconnect_1_utlb_0_ctrl_reg_readdata),        //              .readdata
		.avs_ctrl_reg_waitrequest (mm_interconnect_1_utlb_0_ctrl_reg_waitrequest),     //              .waitrequest
		.clk                      (philosopher_clk_in_clk),                            //         clock.clk
		.reset                    (rst_controller_reset_out_reset),                    //         reset.reset
		.avm_byteenable           (utlb_0_avalon_master_byteenable),                   // avalon_master.byteenable
		.avm_read                 (utlb_0_avalon_master_read),                         //              .read
		.avm_write                (utlb_0_avalon_master_write),                        //              .write
		.avm_writedata            (utlb_0_avalon_master_writedata),                    //              .writedata
		.avm_waitrequest          (utlb_0_avalon_master_waitrequest),                  //              .waitrequest
		.avm_readdata             (utlb_0_avalon_master_readdata),                     //              .readdata
		.avm_address              (utlb_0_avalon_master_address),                      //              .address
		.avs_address              (mm_interconnect_1_utlb_0_avalon_slave_address),     //  avalon_slave.address
		.avs_byteenable           (mm_interconnect_1_utlb_0_avalon_slave_byteenable),  //              .byteenable
		.avs_read                 (mm_interconnect_1_utlb_0_avalon_slave_read),        //              .read
		.avs_write                (mm_interconnect_1_utlb_0_avalon_slave_write),       //              .write
		.avs_writedata            (mm_interconnect_1_utlb_0_avalon_slave_writedata),   //              .writedata
		.avs_waitrequest          (mm_interconnect_1_utlb_0_avalon_slave_waitrequest), //              .waitrequest
		.avs_readdata             (mm_interconnect_1_utlb_0_avalon_slave_readdata),    //              .readdata
		.avs_address_conduit      (),                                                  //       conduit.address
		.fprint_waitrequest       (utlb_0_fprint_waitrequest),                         //        fprint.export
		.fprint_data_address      (utlb_0_fprint_data_address),                        //              .export
		.fprint_writedata         (utlb_0_fprint_writedata),                           //              .export
		.fprint_write             (utlb_0_fprint_write)                                //              .export
	);

	nios_fprint_processor1_0_nios_custom_instr_floating_point_2_0 nios_custom_instr_floating_point_2_0 (
		.s1_dataa     (cpu1_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (cpu1_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (cpu1_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (cpu1_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	nios_fprint_processor1_0_scratchpad_1 scratchpad_1 (
		.clk        (philosopher_clk_in_clk),                       //   clk1.clk
		.address    (mm_interconnect_0_scratchpad_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_scratchpad_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_scratchpad_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_scratchpad_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_scratchpad_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_scratchpad_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_scratchpad_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)            //       .reset_req
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpu1_custom_instruction_master_translator (
		.ci_slave_dataa            (cpu1_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (cpu1_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (cpu1_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (cpu1_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (cpu1_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (cpu1_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (cpu1_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (cpu1_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (cpu1_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (cpu1_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (),                                                                    //                .ipending
		.ci_slave_estatus          (),                                                                    //                .estatus
		.ci_slave_multi_clk        (cpu1_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (cpu1_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (cpu1_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (cpu1_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (cpu1_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (cpu1_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (cpu1_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (cpu1_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (cpu1_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (cpu1_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (cpu1_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (cpu1_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (cpu1_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (cpu1_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (cpu1_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (cpu1_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (cpu1_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (cpu1_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (cpu1_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (cpu1_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (cpu1_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (cpu1_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (cpu1_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (cpu1_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (cpu1_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (cpu1_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (cpu1_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (cpu1_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (cpu1_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (cpu1_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (cpu1_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (cpu1_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (cpu1_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (cpu1_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (cpu1_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (cpu1_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (cpu1_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (cpu1_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (cpu1_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (cpu1_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (cpu1_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (cpu1_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (cpu1_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (cpu1_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	nios_fprint_processor1_0_cpu1_custom_instruction_master_comb_xconnect cpu1_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpu1_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpu1_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpu1_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpu1_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpu1_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpu1_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpu1_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpu1_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpu1_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpu1_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpu1_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpu1_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpu1_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpu1_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpu1_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpu1_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpu1_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpu1_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpu1_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpu1_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpu1_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpu1_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpu1_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpu1_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) cpu1_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (cpu1_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpu1_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpu1_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpu1_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpu1_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpu1_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpu1_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpu1_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpu1_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpu1_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpu1_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpu1_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (cpu1_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpu1_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (cpu1_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (cpu1_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                       // (terminated)
		.ci_master_readrb    (),                                                                       // (terminated)
		.ci_master_writerc   (),                                                                       // (terminated)
		.ci_master_a         (),                                                                       // (terminated)
		.ci_master_b         (),                                                                       // (terminated)
		.ci_master_c         (),                                                                       // (terminated)
		.ci_master_ipending  (),                                                                       // (terminated)
		.ci_master_estatus   (),                                                                       // (terminated)
		.ci_master_clk       (),                                                                       // (terminated)
		.ci_master_clken     (),                                                                       // (terminated)
		.ci_master_reset_req (),                                                                       // (terminated)
		.ci_master_reset     (),                                                                       // (terminated)
		.ci_master_start     (),                                                                       // (terminated)
		.ci_master_done      (1'b0),                                                                   // (terminated)
		.ci_slave_clk        (1'b0),                                                                   // (terminated)
		.ci_slave_clken      (1'b0),                                                                   // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                   // (terminated)
		.ci_slave_reset      (1'b0),                                                                   // (terminated)
		.ci_slave_start      (1'b0),                                                                   // (terminated)
		.ci_slave_done       ()                                                                        // (terminated)
	);

	nios_fprint_processor1_0_cpu1_custom_instruction_master_multi_xconnect cpu1_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (cpu1_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (cpu1_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (cpu1_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (cpu1_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (cpu1_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (cpu1_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (cpu1_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (cpu1_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (cpu1_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (cpu1_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                    //           .ipending
		.ci_slave_estatus     (),                                                                    //           .estatus
		.ci_slave_clk         (cpu1_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (cpu1_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (cpu1_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (cpu1_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (cpu1_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (cpu1_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (cpu1_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (cpu1_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (cpu1_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (cpu1_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (cpu1_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (cpu1_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (cpu1_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (cpu1_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (cpu1_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (cpu1_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (cpu1_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (cpu1_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (cpu1_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (cpu1_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (cpu1_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (cpu1_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (cpu1_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (cpu1_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) cpu1_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (cpu1_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (cpu1_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (cpu1_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (cpu1_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (cpu1_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (cpu1_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (cpu1_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (cpu1_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (cpu1_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (cpu1_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (cpu1_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (cpu1_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (cpu1_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (cpu1_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (cpu1_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (cpu1_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (cpu1_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (cpu1_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (cpu1_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                           // (terminated)
		.ci_master_readrb    (),                                                                           // (terminated)
		.ci_master_writerc   (),                                                                           // (terminated)
		.ci_master_a         (),                                                                           // (terminated)
		.ci_master_b         (),                                                                           // (terminated)
		.ci_master_c         (),                                                                           // (terminated)
		.ci_master_ipending  (),                                                                           // (terminated)
		.ci_master_estatus   ()                                                                            // (terminated)
	);

	nios_fprint_processor1_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                             (philosopher_clk_in_clk),                               //                           clk_clk.clk
		.dma_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // dma_0_reset_reset_bridge_in_reset.reset
		.dma_0_read_master_address               (dma_0_read_master_address),                            //                 dma_0_read_master.address
		.dma_0_read_master_waitrequest           (dma_0_read_master_waitrequest),                        //                                  .waitrequest
		.dma_0_read_master_chipselect            (dma_0_read_master_chipselect),                         //                                  .chipselect
		.dma_0_read_master_read                  (~dma_0_read_master_read),                              //                                  .read
		.dma_0_read_master_readdata              (dma_0_read_master_readdata),                           //                                  .readdata
		.dma_0_read_master_readdatavalid         (dma_0_read_master_readdatavalid),                      //                                  .readdatavalid
		.dma_0_write_master_address              (dma_0_write_master_address),                           //                dma_0_write_master.address
		.dma_0_write_master_waitrequest          (dma_0_write_master_waitrequest),                       //                                  .waitrequest
		.dma_0_write_master_byteenable           (dma_0_write_master_byteenable),                        //                                  .byteenable
		.dma_0_write_master_chipselect           (dma_0_write_master_chipselect),                        //                                  .chipselect
		.dma_0_write_master_write                (~dma_0_write_master_write),                            //                                  .write
		.dma_0_write_master_writedata            (dma_0_write_master_writedata),                         //                                  .writedata
		.utlb_0_avalon_master_address            (utlb_0_avalon_master_address),                         //              utlb_0_avalon_master.address
		.utlb_0_avalon_master_waitrequest        (utlb_0_avalon_master_waitrequest),                     //                                  .waitrequest
		.utlb_0_avalon_master_byteenable         (utlb_0_avalon_master_byteenable),                      //                                  .byteenable
		.utlb_0_avalon_master_read               (utlb_0_avalon_master_read),                            //                                  .read
		.utlb_0_avalon_master_readdata           (utlb_0_avalon_master_readdata),                        //                                  .readdata
		.utlb_0_avalon_master_write              (utlb_0_avalon_master_write),                           //                                  .write
		.utlb_0_avalon_master_writedata          (utlb_0_avalon_master_writedata),                       //                                  .writedata
		.out_system_bridge_s0_address            (mm_interconnect_0_out_system_bridge_s0_address),       //              out_system_bridge_s0.address
		.out_system_bridge_s0_write              (mm_interconnect_0_out_system_bridge_s0_write),         //                                  .write
		.out_system_bridge_s0_read               (mm_interconnect_0_out_system_bridge_s0_read),          //                                  .read
		.out_system_bridge_s0_readdata           (mm_interconnect_0_out_system_bridge_s0_readdata),      //                                  .readdata
		.out_system_bridge_s0_writedata          (mm_interconnect_0_out_system_bridge_s0_writedata),     //                                  .writedata
		.out_system_bridge_s0_burstcount         (mm_interconnect_0_out_system_bridge_s0_burstcount),    //                                  .burstcount
		.out_system_bridge_s0_byteenable         (mm_interconnect_0_out_system_bridge_s0_byteenable),    //                                  .byteenable
		.out_system_bridge_s0_readdatavalid      (mm_interconnect_0_out_system_bridge_s0_readdatavalid), //                                  .readdatavalid
		.out_system_bridge_s0_waitrequest        (mm_interconnect_0_out_system_bridge_s0_waitrequest),   //                                  .waitrequest
		.out_system_bridge_s0_debugaccess        (mm_interconnect_0_out_system_bridge_s0_debugaccess),   //                                  .debugaccess
		.scratchpad_0_s1_address                 (mm_interconnect_0_scratchpad_0_s1_address),            //                   scratchpad_0_s1.address
		.scratchpad_0_s1_write                   (mm_interconnect_0_scratchpad_0_s1_write),              //                                  .write
		.scratchpad_0_s1_readdata                (mm_interconnect_0_scratchpad_0_s1_readdata),           //                                  .readdata
		.scratchpad_0_s1_writedata               (mm_interconnect_0_scratchpad_0_s1_writedata),          //                                  .writedata
		.scratchpad_0_s1_byteenable              (mm_interconnect_0_scratchpad_0_s1_byteenable),         //                                  .byteenable
		.scratchpad_0_s1_chipselect              (mm_interconnect_0_scratchpad_0_s1_chipselect),         //                                  .chipselect
		.scratchpad_0_s1_clken                   (mm_interconnect_0_scratchpad_0_s1_clken),              //                                  .clken
		.scratchpad_1_s1_address                 (mm_interconnect_0_scratchpad_1_s1_address),            //                   scratchpad_1_s1.address
		.scratchpad_1_s1_write                   (mm_interconnect_0_scratchpad_1_s1_write),              //                                  .write
		.scratchpad_1_s1_readdata                (mm_interconnect_0_scratchpad_1_s1_readdata),           //                                  .readdata
		.scratchpad_1_s1_writedata               (mm_interconnect_0_scratchpad_1_s1_writedata),          //                                  .writedata
		.scratchpad_1_s1_byteenable              (mm_interconnect_0_scratchpad_1_s1_byteenable),         //                                  .byteenable
		.scratchpad_1_s1_chipselect              (mm_interconnect_0_scratchpad_1_s1_chipselect),         //                                  .chipselect
		.scratchpad_1_s1_clken                   (mm_interconnect_0_scratchpad_1_s1_clken)               //                                  .clken
	);

	nios_fprint_processor1_0_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                              (philosopher_clk_in_clk),                                     //                            clk_clk.clk
		.cpu1_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                             // cpu1_reset_n_reset_bridge_in_reset.reset
		.cpu1_data_master_address                 (cpu1_data_master_address),                                   //                   cpu1_data_master.address
		.cpu1_data_master_waitrequest             (cpu1_data_master_waitrequest),                               //                                   .waitrequest
		.cpu1_data_master_byteenable              (cpu1_data_master_byteenable),                                //                                   .byteenable
		.cpu1_data_master_read                    (cpu1_data_master_read),                                      //                                   .read
		.cpu1_data_master_readdata                (cpu1_data_master_readdata),                                  //                                   .readdata
		.cpu1_data_master_write                   (cpu1_data_master_write),                                     //                                   .write
		.cpu1_data_master_writedata               (cpu1_data_master_writedata),                                 //                                   .writedata
		.cpu1_data_master_debugaccess             (cpu1_data_master_debugaccess),                               //                                   .debugaccess
		.cpu1_instruction_master_address          (cpu1_instruction_master_address),                            //            cpu1_instruction_master.address
		.cpu1_instruction_master_waitrequest      (cpu1_instruction_master_waitrequest),                        //                                   .waitrequest
		.cpu1_instruction_master_read             (cpu1_instruction_master_read),                               //                                   .read
		.cpu1_instruction_master_readdata         (cpu1_instruction_master_readdata),                           //                                   .readdata
		.cpu1_instruction_master_readdatavalid    (cpu1_instruction_master_readdatavalid),                      //                                   .readdatavalid
		.cpu1_jtag_debug_module_address           (mm_interconnect_1_cpu1_jtag_debug_module_address),           //             cpu1_jtag_debug_module.address
		.cpu1_jtag_debug_module_write             (mm_interconnect_1_cpu1_jtag_debug_module_write),             //                                   .write
		.cpu1_jtag_debug_module_read              (mm_interconnect_1_cpu1_jtag_debug_module_read),              //                                   .read
		.cpu1_jtag_debug_module_readdata          (mm_interconnect_1_cpu1_jtag_debug_module_readdata),          //                                   .readdata
		.cpu1_jtag_debug_module_writedata         (mm_interconnect_1_cpu1_jtag_debug_module_writedata),         //                                   .writedata
		.cpu1_jtag_debug_module_byteenable        (mm_interconnect_1_cpu1_jtag_debug_module_byteenable),        //                                   .byteenable
		.cpu1_jtag_debug_module_waitrequest       (mm_interconnect_1_cpu1_jtag_debug_module_waitrequest),       //                                   .waitrequest
		.cpu1_jtag_debug_module_debugaccess       (mm_interconnect_1_cpu1_jtag_debug_module_debugaccess),       //                                   .debugaccess
		.Fingerprint_0_avalon_slave_0_address     (mm_interconnect_1_fingerprint_0_avalon_slave_0_address),     //       Fingerprint_0_avalon_slave_0.address
		.Fingerprint_0_avalon_slave_0_write       (mm_interconnect_1_fingerprint_0_avalon_slave_0_write),       //                                   .write
		.Fingerprint_0_avalon_slave_0_read        (mm_interconnect_1_fingerprint_0_avalon_slave_0_read),        //                                   .read
		.Fingerprint_0_avalon_slave_0_readdata    (mm_interconnect_1_fingerprint_0_avalon_slave_0_readdata),    //                                   .readdata
		.Fingerprint_0_avalon_slave_0_writedata   (mm_interconnect_1_fingerprint_0_avalon_slave_0_writedata),   //                                   .writedata
		.Fingerprint_0_avalon_slave_0_waitrequest (mm_interconnect_1_fingerprint_0_avalon_slave_0_waitrequest), //                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_address      (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),      //        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),        //                                   .write
		.jtag_uart_avalon_jtag_slave_read         (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),         //                                   .read
		.jtag_uart_avalon_jtag_slave_readdata     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),     //                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),    //                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),  //                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),   //                                   .chipselect
		.timer_s1_address                         (mm_interconnect_1_timer_s1_address),                         //                           timer_s1.address
		.timer_s1_write                           (mm_interconnect_1_timer_s1_write),                           //                                   .write
		.timer_s1_readdata                        (mm_interconnect_1_timer_s1_readdata),                        //                                   .readdata
		.timer_s1_writedata                       (mm_interconnect_1_timer_s1_writedata),                       //                                   .writedata
		.timer_s1_chipselect                      (mm_interconnect_1_timer_s1_chipselect),                      //                                   .chipselect
		.timestamp_s1_address                     (mm_interconnect_1_timestamp_s1_address),                     //                       timestamp_s1.address
		.timestamp_s1_write                       (mm_interconnect_1_timestamp_s1_write),                       //                                   .write
		.timestamp_s1_readdata                    (mm_interconnect_1_timestamp_s1_readdata),                    //                                   .readdata
		.timestamp_s1_writedata                   (mm_interconnect_1_timestamp_s1_writedata),                   //                                   .writedata
		.timestamp_s1_chipselect                  (mm_interconnect_1_timestamp_s1_chipselect),                  //                                   .chipselect
		.utlb_0_avalon_slave_address              (mm_interconnect_1_utlb_0_avalon_slave_address),              //                utlb_0_avalon_slave.address
		.utlb_0_avalon_slave_write                (mm_interconnect_1_utlb_0_avalon_slave_write),                //                                   .write
		.utlb_0_avalon_slave_read                 (mm_interconnect_1_utlb_0_avalon_slave_read),                 //                                   .read
		.utlb_0_avalon_slave_readdata             (mm_interconnect_1_utlb_0_avalon_slave_readdata),             //                                   .readdata
		.utlb_0_avalon_slave_writedata            (mm_interconnect_1_utlb_0_avalon_slave_writedata),            //                                   .writedata
		.utlb_0_avalon_slave_byteenable           (mm_interconnect_1_utlb_0_avalon_slave_byteenable),           //                                   .byteenable
		.utlb_0_avalon_slave_waitrequest          (mm_interconnect_1_utlb_0_avalon_slave_waitrequest),          //                                   .waitrequest
		.utlb_0_ctrl_reg_address                  (mm_interconnect_1_utlb_0_ctrl_reg_address),                  //                    utlb_0_ctrl_reg.address
		.utlb_0_ctrl_reg_write                    (mm_interconnect_1_utlb_0_ctrl_reg_write),                    //                                   .write
		.utlb_0_ctrl_reg_read                     (mm_interconnect_1_utlb_0_ctrl_reg_read),                     //                                   .read
		.utlb_0_ctrl_reg_readdata                 (mm_interconnect_1_utlb_0_ctrl_reg_readdata),                 //                                   .readdata
		.utlb_0_ctrl_reg_writedata                (mm_interconnect_1_utlb_0_ctrl_reg_writedata),                //                                   .writedata
		.utlb_0_ctrl_reg_waitrequest              (mm_interconnect_1_utlb_0_ctrl_reg_waitrequest)               //                                   .waitrequest
	);

	nios_fprint_processor1_0_irq_mapper irq_mapper (
		.clk           (philosopher_clk_in_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu1_d_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (philosopher_clk_in_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
