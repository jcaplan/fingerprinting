library verilog;
use verilog.vl_types.all;
entity tb_comp_registers is
end tb_comp_registers;
