library verilog;
use verilog.vl_types.all;
entity tb_comparator is
end tb_comparator;
