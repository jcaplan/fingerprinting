library verilog;
use verilog.vl_types.all;
entity tb_csr_registers is
end tb_csr_registers;
