library verilog;
use verilog.vl_types.all;
entity tb_fprint_registers is
end tb_fprint_registers;
