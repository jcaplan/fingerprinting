`include "crc_defines.v"
module csr_decode(
	input										clk,
	input										reset,
	input 	[(`COMPARATOR_ADDRESS_WIDTH-1):0]	fprint_address,
	input 	[(`NIOS_DATA_WIDTH-1):0]			fprint_writedata,
	



);


//we need the index to do this properly... have to go start in the registers file...

endmodule
