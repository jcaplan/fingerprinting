// nios_fprint_processorM_0.v

// Generated using ACDS version 13.1 162 at 2016.01.16.18:27:46

`timescale 1 ps / 1 ps
module nios_fprint_processorM_0 (
		input  wire        philosopher_clk_in_clk,                //             philosopher_clk_in.clk
		input  wire        outgoing_master_waitrequest,           //                outgoing_master.waitrequest
		input  wire [31:0] outgoing_master_readdata,              //                               .readdata
		input  wire        outgoing_master_readdatavalid,         //                               .readdatavalid
		output wire [0:0]  outgoing_master_burstcount,            //                               .burstcount
		output wire [31:0] outgoing_master_writedata,             //                               .writedata
		output wire [26:0] outgoing_master_address,               //                               .address
		output wire        outgoing_master_write,                 //                               .write
		output wire        outgoing_master_read,                  //                               .read
		output wire [3:0]  outgoing_master_byteenable,            //                               .byteenable
		output wire        outgoing_master_debugaccess,           //                               .debugaccess
		input  wire        button_pio_external_connection_export, // button_pio_external_connection.export
		output wire        cpu0_jtag_debug_module_reset_reset,    //   cpu0_jtag_debug_module_reset.reset
		input  wire        reset_reset_n,                         //                          reset.reset_n
		input  wire        fprint_irq_0_irq_export,               //               fprint_irq_0_irq.export
		input  wire [7:0]  cpu_irq_0_s0_address,                  //                   cpu_irq_0_s0.address
		input  wire        cpu_irq_0_s0_write,                    //                               .write
		input  wire [31:0] cpu_irq_0_s0_writedata,                //                               .writedata
		input  wire [7:0]  reset_monitor_0_s0_address,            //             reset_monitor_0_s0.address
		input  wire        reset_monitor_0_s0_read,               //                               .read
		output wire [31:0] reset_monitor_0_s0_readdata,           //                               .readdata
		input  wire        reset_monitor_0_s0_write,              //                               .write
		input  wire [31:0] reset_monitor_0_s0_writedata,          //                               .writedata
		output wire        reset_monitor_0_s0_waitrequest,        //                               .waitrequest
		input  wire [3:0]  dma_0_irq_receiver_irq_irq             //         dma_0_irq_receiver_irq.irq
	);

	wire  [31:0] cpum_custom_instruction_master_result;                                      // cpuM_custom_instruction_master_translator:ci_slave_result -> cpuM:E_ci_combo_result
	wire   [7:0] cpum_custom_instruction_master_multi_n;                                     // cpuM:A_ci_multi_n -> cpuM_custom_instruction_master_translator:ci_slave_multi_n
	wire         cpum_custom_instruction_master_writerc;                                     // cpuM:E_ci_combo_writerc -> cpuM_custom_instruction_master_translator:ci_slave_writerc
	wire  [31:0] cpum_custom_instruction_master_multi_result;                                // cpuM_custom_instruction_master_translator:ci_slave_multi_result -> cpuM:A_ci_multi_result
	wire  [31:0] cpum_custom_instruction_master_multi_dataa;                                 // cpuM:A_ci_multi_dataa -> cpuM_custom_instruction_master_translator:ci_slave_multi_dataa
	wire  [31:0] cpum_custom_instruction_master_dataa;                                       // cpuM:E_ci_combo_dataa -> cpuM_custom_instruction_master_translator:ci_slave_dataa
	wire  [31:0] cpum_custom_instruction_master_multi_datab;                                 // cpuM:A_ci_multi_datab -> cpuM_custom_instruction_master_translator:ci_slave_multi_datab
	wire         cpum_custom_instruction_master_readra;                                      // cpuM:E_ci_combo_readra -> cpuM_custom_instruction_master_translator:ci_slave_readra
	wire         cpum_custom_instruction_master_reset;                                       // cpuM:A_ci_multi_reset -> cpuM_custom_instruction_master_translator:ci_slave_multi_reset
	wire  [31:0] cpum_custom_instruction_master_datab;                                       // cpuM:E_ci_combo_datab -> cpuM_custom_instruction_master_translator:ci_slave_datab
	wire         cpum_custom_instruction_master_readrb;                                      // cpuM:E_ci_combo_readrb -> cpuM_custom_instruction_master_translator:ci_slave_readrb
	wire         cpum_custom_instruction_master_multi_readra;                                // cpuM:A_ci_multi_readra -> cpuM_custom_instruction_master_translator:ci_slave_multi_readra
	wire         cpum_custom_instruction_master_multi_readrb;                                // cpuM:A_ci_multi_readrb -> cpuM_custom_instruction_master_translator:ci_slave_multi_readrb
	wire   [4:0] cpum_custom_instruction_master_b;                                           // cpuM:E_ci_combo_b -> cpuM_custom_instruction_master_translator:ci_slave_b
	wire   [4:0] cpum_custom_instruction_master_c;                                           // cpuM:E_ci_combo_c -> cpuM_custom_instruction_master_translator:ci_slave_c
	wire         cpum_custom_instruction_master_clk_en;                                      // cpuM:A_ci_multi_clk_en -> cpuM_custom_instruction_master_translator:ci_slave_multi_clken
	wire         cpum_custom_instruction_master_done;                                        // cpuM_custom_instruction_master_translator:ci_slave_multi_done -> cpuM:A_ci_multi_done
	wire   [4:0] cpum_custom_instruction_master_a;                                           // cpuM:E_ci_combo_a -> cpuM_custom_instruction_master_translator:ci_slave_a
	wire   [7:0] cpum_custom_instruction_master_n;                                           // cpuM:E_ci_combo_n -> cpuM_custom_instruction_master_translator:ci_slave_n
	wire         cpum_custom_instruction_master_multi_writerc;                               // cpuM:A_ci_multi_writerc -> cpuM_custom_instruction_master_translator:ci_slave_multi_writerc
	wire         cpum_custom_instruction_master_clk;                                         // cpuM:A_ci_multi_clock -> cpuM_custom_instruction_master_translator:ci_slave_multi_clk
	wire         cpum_custom_instruction_master_reset_req;                                   // cpuM:A_ci_multi_reset_req -> cpuM_custom_instruction_master_translator:ci_slave_multi_reset_req
	wire   [4:0] cpum_custom_instruction_master_multi_c;                                     // cpuM:A_ci_multi_c -> cpuM_custom_instruction_master_translator:ci_slave_multi_c
	wire   [4:0] cpum_custom_instruction_master_multi_b;                                     // cpuM:A_ci_multi_b -> cpuM_custom_instruction_master_translator:ci_slave_multi_b
	wire   [4:0] cpum_custom_instruction_master_multi_a;                                     // cpuM:A_ci_multi_a -> cpuM_custom_instruction_master_translator:ci_slave_multi_a
	wire         cpum_custom_instruction_master_start;                                       // cpuM:A_ci_multi_start -> cpuM_custom_instruction_master_translator:ci_slave_multi_start
	wire  [31:0] cpum_custom_instruction_master_translator_comb_ci_master_result;            // cpuM_custom_instruction_master_comb_xconnect:ci_slave_result -> cpuM_custom_instruction_master_translator:comb_ci_master_result
	wire   [4:0] cpum_custom_instruction_master_translator_comb_ci_master_b;                 // cpuM_custom_instruction_master_translator:comb_ci_master_b -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_b
	wire   [4:0] cpum_custom_instruction_master_translator_comb_ci_master_c;                 // cpuM_custom_instruction_master_translator:comb_ci_master_c -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_c
	wire  [31:0] cpum_custom_instruction_master_translator_comb_ci_master_dataa;             // cpuM_custom_instruction_master_translator:comb_ci_master_dataa -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_dataa
	wire   [4:0] cpum_custom_instruction_master_translator_comb_ci_master_a;                 // cpuM_custom_instruction_master_translator:comb_ci_master_a -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_a
	wire         cpum_custom_instruction_master_translator_comb_ci_master_readra;            // cpuM_custom_instruction_master_translator:comb_ci_master_readra -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_readra
	wire   [7:0] cpum_custom_instruction_master_translator_comb_ci_master_n;                 // cpuM_custom_instruction_master_translator:comb_ci_master_n -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_n
	wire         cpum_custom_instruction_master_translator_comb_ci_master_writerc;           // cpuM_custom_instruction_master_translator:comb_ci_master_writerc -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_writerc
	wire  [31:0] cpum_custom_instruction_master_translator_comb_ci_master_datab;             // cpuM_custom_instruction_master_translator:comb_ci_master_datab -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_datab
	wire  [31:0] cpum_custom_instruction_master_translator_comb_ci_master_ipending;          // cpuM_custom_instruction_master_translator:comb_ci_master_ipending -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_ipending
	wire         cpum_custom_instruction_master_translator_comb_ci_master_readrb;            // cpuM_custom_instruction_master_translator:comb_ci_master_readrb -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_readrb
	wire         cpum_custom_instruction_master_translator_comb_ci_master_estatus;           // cpuM_custom_instruction_master_translator:comb_ci_master_estatus -> cpuM_custom_instruction_master_comb_xconnect:ci_slave_estatus
	wire  [31:0] cpum_custom_instruction_master_comb_xconnect_ci_master0_result;             // cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_result -> cpuM_custom_instruction_master_comb_xconnect:ci_master0_result
	wire   [4:0] cpum_custom_instruction_master_comb_xconnect_ci_master0_b;                  // cpuM_custom_instruction_master_comb_xconnect:ci_master0_b -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_b
	wire   [4:0] cpum_custom_instruction_master_comb_xconnect_ci_master0_c;                  // cpuM_custom_instruction_master_comb_xconnect:ci_master0_c -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_c
	wire  [31:0] cpum_custom_instruction_master_comb_xconnect_ci_master0_dataa;              // cpuM_custom_instruction_master_comb_xconnect:ci_master0_dataa -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_dataa
	wire   [4:0] cpum_custom_instruction_master_comb_xconnect_ci_master0_a;                  // cpuM_custom_instruction_master_comb_xconnect:ci_master0_a -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_a
	wire         cpum_custom_instruction_master_comb_xconnect_ci_master0_readra;             // cpuM_custom_instruction_master_comb_xconnect:ci_master0_readra -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_readra
	wire   [7:0] cpum_custom_instruction_master_comb_xconnect_ci_master0_n;                  // cpuM_custom_instruction_master_comb_xconnect:ci_master0_n -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_n
	wire         cpum_custom_instruction_master_comb_xconnect_ci_master0_writerc;            // cpuM_custom_instruction_master_comb_xconnect:ci_master0_writerc -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_writerc
	wire  [31:0] cpum_custom_instruction_master_comb_xconnect_ci_master0_datab;              // cpuM_custom_instruction_master_comb_xconnect:ci_master0_datab -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_datab
	wire  [31:0] cpum_custom_instruction_master_comb_xconnect_ci_master0_ipending;           // cpuM_custom_instruction_master_comb_xconnect:ci_master0_ipending -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_ipending
	wire         cpum_custom_instruction_master_comb_xconnect_ci_master0_readrb;             // cpuM_custom_instruction_master_comb_xconnect:ci_master0_readrb -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_readrb
	wire         cpum_custom_instruction_master_comb_xconnect_ci_master0_estatus;            // cpuM_custom_instruction_master_comb_xconnect:ci_master0_estatus -> cpuM_custom_instruction_master_comb_slave_translator0:ci_slave_estatus
	wire  [31:0] cpum_custom_instruction_master_comb_slave_translator0_ci_master_result;     // nios_custom_instr_floating_point_2_0:s1_result -> cpuM_custom_instruction_master_comb_slave_translator0:ci_master_result
	wire  [31:0] cpum_custom_instruction_master_comb_slave_translator0_ci_master_dataa;      // cpuM_custom_instruction_master_comb_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s1_dataa
	wire   [3:0] cpum_custom_instruction_master_comb_slave_translator0_ci_master_n;          // cpuM_custom_instruction_master_comb_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s1_n
	wire  [31:0] cpum_custom_instruction_master_comb_slave_translator0_ci_master_datab;      // cpuM_custom_instruction_master_comb_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s1_datab
	wire  [31:0] cpum_custom_instruction_master_translator_multi_ci_master_result;           // cpuM_custom_instruction_master_multi_xconnect:ci_slave_result -> cpuM_custom_instruction_master_translator:multi_ci_master_result
	wire   [4:0] cpum_custom_instruction_master_translator_multi_ci_master_b;                // cpuM_custom_instruction_master_translator:multi_ci_master_b -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_b
	wire   [4:0] cpum_custom_instruction_master_translator_multi_ci_master_c;                // cpuM_custom_instruction_master_translator:multi_ci_master_c -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_c
	wire   [4:0] cpum_custom_instruction_master_translator_multi_ci_master_a;                // cpuM_custom_instruction_master_translator:multi_ci_master_a -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_a
	wire         cpum_custom_instruction_master_translator_multi_ci_master_clk_en;           // cpuM_custom_instruction_master_translator:multi_ci_master_clken -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_clken
	wire         cpum_custom_instruction_master_translator_multi_ci_master_done;             // cpuM_custom_instruction_master_multi_xconnect:ci_slave_done -> cpuM_custom_instruction_master_translator:multi_ci_master_done
	wire   [7:0] cpum_custom_instruction_master_translator_multi_ci_master_n;                // cpuM_custom_instruction_master_translator:multi_ci_master_n -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_n
	wire         cpum_custom_instruction_master_translator_multi_ci_master_writerc;          // cpuM_custom_instruction_master_translator:multi_ci_master_writerc -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_writerc
	wire         cpum_custom_instruction_master_translator_multi_ci_master_clk;              // cpuM_custom_instruction_master_translator:multi_ci_master_clk -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_clk
	wire         cpum_custom_instruction_master_translator_multi_ci_master_reset_req;        // cpuM_custom_instruction_master_translator:multi_ci_master_reset_req -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_reset_req
	wire         cpum_custom_instruction_master_translator_multi_ci_master_start;            // cpuM_custom_instruction_master_translator:multi_ci_master_start -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_start
	wire  [31:0] cpum_custom_instruction_master_translator_multi_ci_master_dataa;            // cpuM_custom_instruction_master_translator:multi_ci_master_dataa -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_dataa
	wire         cpum_custom_instruction_master_translator_multi_ci_master_readra;           // cpuM_custom_instruction_master_translator:multi_ci_master_readra -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_readra
	wire         cpum_custom_instruction_master_translator_multi_ci_master_reset;            // cpuM_custom_instruction_master_translator:multi_ci_master_reset -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_reset
	wire  [31:0] cpum_custom_instruction_master_translator_multi_ci_master_datab;            // cpuM_custom_instruction_master_translator:multi_ci_master_datab -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_datab
	wire         cpum_custom_instruction_master_translator_multi_ci_master_readrb;           // cpuM_custom_instruction_master_translator:multi_ci_master_readrb -> cpuM_custom_instruction_master_multi_xconnect:ci_slave_readrb
	wire  [31:0] cpum_custom_instruction_master_multi_xconnect_ci_master0_result;            // cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_result -> cpuM_custom_instruction_master_multi_xconnect:ci_master0_result
	wire   [4:0] cpum_custom_instruction_master_multi_xconnect_ci_master0_b;                 // cpuM_custom_instruction_master_multi_xconnect:ci_master0_b -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_b
	wire   [4:0] cpum_custom_instruction_master_multi_xconnect_ci_master0_c;                 // cpuM_custom_instruction_master_multi_xconnect:ci_master0_c -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_c
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_done;              // cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_done -> cpuM_custom_instruction_master_multi_xconnect:ci_master0_done
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_clk_en;            // cpuM_custom_instruction_master_multi_xconnect:ci_master0_clken -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_clken
	wire   [4:0] cpum_custom_instruction_master_multi_xconnect_ci_master0_a;                 // cpuM_custom_instruction_master_multi_xconnect:ci_master0_a -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_a
	wire   [7:0] cpum_custom_instruction_master_multi_xconnect_ci_master0_n;                 // cpuM_custom_instruction_master_multi_xconnect:ci_master0_n -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_n
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_writerc;           // cpuM_custom_instruction_master_multi_xconnect:ci_master0_writerc -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_writerc
	wire  [31:0] cpum_custom_instruction_master_multi_xconnect_ci_master0_ipending;          // cpuM_custom_instruction_master_multi_xconnect:ci_master0_ipending -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_ipending
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_clk;               // cpuM_custom_instruction_master_multi_xconnect:ci_master0_clk -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_clk
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_reset_req;         // cpuM_custom_instruction_master_multi_xconnect:ci_master0_reset_req -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_reset_req
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_start;             // cpuM_custom_instruction_master_multi_xconnect:ci_master0_start -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_start
	wire  [31:0] cpum_custom_instruction_master_multi_xconnect_ci_master0_dataa;             // cpuM_custom_instruction_master_multi_xconnect:ci_master0_dataa -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_dataa
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_readra;            // cpuM_custom_instruction_master_multi_xconnect:ci_master0_readra -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_readra
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_reset;             // cpuM_custom_instruction_master_multi_xconnect:ci_master0_reset -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_reset
	wire  [31:0] cpum_custom_instruction_master_multi_xconnect_ci_master0_datab;             // cpuM_custom_instruction_master_multi_xconnect:ci_master0_datab -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_datab
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_readrb;            // cpuM_custom_instruction_master_multi_xconnect:ci_master0_readrb -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_readrb
	wire         cpum_custom_instruction_master_multi_xconnect_ci_master0_estatus;           // cpuM_custom_instruction_master_multi_xconnect:ci_master0_estatus -> cpuM_custom_instruction_master_multi_slave_translator0:ci_slave_estatus
	wire  [31:0] cpum_custom_instruction_master_multi_slave_translator0_ci_master_result;    // nios_custom_instr_floating_point_2_0:s2_result -> cpuM_custom_instruction_master_multi_slave_translator0:ci_master_result
	wire         cpum_custom_instruction_master_multi_slave_translator0_ci_master_start;     // cpuM_custom_instruction_master_multi_slave_translator0:ci_master_start -> nios_custom_instr_floating_point_2_0:s2_start
	wire  [31:0] cpum_custom_instruction_master_multi_slave_translator0_ci_master_dataa;     // cpuM_custom_instruction_master_multi_slave_translator0:ci_master_dataa -> nios_custom_instr_floating_point_2_0:s2_dataa
	wire         cpum_custom_instruction_master_multi_slave_translator0_ci_master_done;      // nios_custom_instr_floating_point_2_0:s2_done -> cpuM_custom_instruction_master_multi_slave_translator0:ci_master_done
	wire         cpum_custom_instruction_master_multi_slave_translator0_ci_master_clk_en;    // cpuM_custom_instruction_master_multi_slave_translator0:ci_master_clken -> nios_custom_instr_floating_point_2_0:s2_clk_en
	wire   [2:0] cpum_custom_instruction_master_multi_slave_translator0_ci_master_n;         // cpuM_custom_instruction_master_multi_slave_translator0:ci_master_n -> nios_custom_instr_floating_point_2_0:s2_n
	wire         cpum_custom_instruction_master_multi_slave_translator0_ci_master_reset;     // cpuM_custom_instruction_master_multi_slave_translator0:ci_master_reset -> nios_custom_instr_floating_point_2_0:s2_reset
	wire  [31:0] cpum_custom_instruction_master_multi_slave_translator0_ci_master_datab;     // cpuM_custom_instruction_master_multi_slave_translator0:ci_master_datab -> nios_custom_instr_floating_point_2_0:s2_datab
	wire         cpum_custom_instruction_master_multi_slave_translator0_ci_master_clk;       // cpuM_custom_instruction_master_multi_slave_translator0:ci_master_clk -> nios_custom_instr_floating_point_2_0:s2_clk
	wire         cpum_custom_instruction_master_multi_slave_translator0_ci_master_reset_req; // cpuM_custom_instruction_master_multi_slave_translator0:ci_master_reset_req -> nios_custom_instr_floating_point_2_0:s2_reset_req
	wire         cpum_instruction_master_waitrequest;                                        // mm_interconnect_0:cpuM_instruction_master_waitrequest -> cpuM:i_waitrequest
	wire  [27:0] cpum_instruction_master_address;                                            // cpuM:i_address -> mm_interconnect_0:cpuM_instruction_master_address
	wire         cpum_instruction_master_read;                                               // cpuM:i_read -> mm_interconnect_0:cpuM_instruction_master_read
	wire  [31:0] cpum_instruction_master_readdata;                                           // mm_interconnect_0:cpuM_instruction_master_readdata -> cpuM:i_readdata
	wire         cpum_instruction_master_readdatavalid;                                      // mm_interconnect_0:cpuM_instruction_master_readdatavalid -> cpuM:i_readdatavalid
	wire  [31:0] mm_interconnect_0_scratchpad_s1_writedata;                                  // mm_interconnect_0:scratchpad_s1_writedata -> scratchpad:writedata
	wire  [11:0] mm_interconnect_0_scratchpad_s1_address;                                    // mm_interconnect_0:scratchpad_s1_address -> scratchpad:address
	wire         mm_interconnect_0_scratchpad_s1_chipselect;                                 // mm_interconnect_0:scratchpad_s1_chipselect -> scratchpad:chipselect
	wire         mm_interconnect_0_scratchpad_s1_clken;                                      // mm_interconnect_0:scratchpad_s1_clken -> scratchpad:clken
	wire         mm_interconnect_0_scratchpad_s1_write;                                      // mm_interconnect_0:scratchpad_s1_write -> scratchpad:write
	wire  [31:0] mm_interconnect_0_scratchpad_s1_readdata;                                   // scratchpad:readdata -> mm_interconnect_0:scratchpad_s1_readdata
	wire   [3:0] mm_interconnect_0_scratchpad_s1_byteenable;                                 // mm_interconnect_0:scratchpad_s1_byteenable -> scratchpad:byteenable
	wire         cpum_data_master_waitrequest;                                               // mm_interconnect_0:cpuM_data_master_waitrequest -> cpuM:d_waitrequest
	wire  [31:0] cpum_data_master_writedata;                                                 // cpuM:d_writedata -> mm_interconnect_0:cpuM_data_master_writedata
	wire  [27:0] cpum_data_master_address;                                                   // cpuM:d_address -> mm_interconnect_0:cpuM_data_master_address
	wire         cpum_data_master_write;                                                     // cpuM:d_write -> mm_interconnect_0:cpuM_data_master_write
	wire         cpum_data_master_read;                                                      // cpuM:d_read -> mm_interconnect_0:cpuM_data_master_read
	wire  [31:0] cpum_data_master_readdata;                                                  // mm_interconnect_0:cpuM_data_master_readdata -> cpuM:d_readdata
	wire         cpum_data_master_debugaccess;                                               // cpuM:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpuM_data_master_debugaccess
	wire   [3:0] cpum_data_master_byteenable;                                                // cpuM:d_byteenable -> mm_interconnect_0:cpuM_data_master_byteenable
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_cpum_jtag_debug_module_waitrequest;                       // cpuM:jtag_debug_module_waitrequest -> mm_interconnect_0:cpuM_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpum_jtag_debug_module_writedata;                         // mm_interconnect_0:cpuM_jtag_debug_module_writedata -> cpuM:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpum_jtag_debug_module_address;                           // mm_interconnect_0:cpuM_jtag_debug_module_address -> cpuM:jtag_debug_module_address
	wire         mm_interconnect_0_cpum_jtag_debug_module_write;                             // mm_interconnect_0:cpuM_jtag_debug_module_write -> cpuM:jtag_debug_module_write
	wire         mm_interconnect_0_cpum_jtag_debug_module_read;                              // mm_interconnect_0:cpuM_jtag_debug_module_read -> cpuM:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpum_jtag_debug_module_readdata;                          // cpuM:jtag_debug_module_readdata -> mm_interconnect_0:cpuM_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpum_jtag_debug_module_debugaccess;                       // mm_interconnect_0:cpuM_jtag_debug_module_debugaccess -> cpuM:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpum_jtag_debug_module_byteenable;                        // mm_interconnect_0:cpuM_jtag_debug_module_byteenable -> cpuM:jtag_debug_module_byteenable
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                       // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                         // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_chipselect;                                      // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire         mm_interconnect_0_timer_s1_write;                                           // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                        // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire  [15:0] mm_interconnect_0_timestamp_s1_writedata;                                   // mm_interconnect_0:timestamp_s1_writedata -> timestamp:writedata
	wire   [3:0] mm_interconnect_0_timestamp_s1_address;                                     // mm_interconnect_0:timestamp_s1_address -> timestamp:address
	wire         mm_interconnect_0_timestamp_s1_chipselect;                                  // mm_interconnect_0:timestamp_s1_chipselect -> timestamp:chipselect
	wire         mm_interconnect_0_timestamp_s1_write;                                       // mm_interconnect_0:timestamp_s1_write -> timestamp:write_n
	wire  [15:0] mm_interconnect_0_timestamp_s1_readdata;                                    // timestamp:readdata -> mm_interconnect_0:timestamp_s1_readdata
	wire         mm_interconnect_0_out_system_bridge_s0_waitrequest;                         // out_system_bridge:s0_waitrequest -> mm_interconnect_0:out_system_bridge_s0_waitrequest
	wire   [0:0] mm_interconnect_0_out_system_bridge_s0_burstcount;                          // mm_interconnect_0:out_system_bridge_s0_burstcount -> out_system_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_writedata;                           // mm_interconnect_0:out_system_bridge_s0_writedata -> out_system_bridge:s0_writedata
	wire  [26:0] mm_interconnect_0_out_system_bridge_s0_address;                             // mm_interconnect_0:out_system_bridge_s0_address -> out_system_bridge:s0_address
	wire         mm_interconnect_0_out_system_bridge_s0_write;                               // mm_interconnect_0:out_system_bridge_s0_write -> out_system_bridge:s0_write
	wire         mm_interconnect_0_out_system_bridge_s0_read;                                // mm_interconnect_0:out_system_bridge_s0_read -> out_system_bridge:s0_read
	wire  [31:0] mm_interconnect_0_out_system_bridge_s0_readdata;                            // out_system_bridge:s0_readdata -> mm_interconnect_0:out_system_bridge_s0_readdata
	wire         mm_interconnect_0_out_system_bridge_s0_debugaccess;                         // mm_interconnect_0:out_system_bridge_s0_debugaccess -> out_system_bridge:s0_debugaccess
	wire         mm_interconnect_0_out_system_bridge_s0_readdatavalid;                       // out_system_bridge:s0_readdatavalid -> mm_interconnect_0:out_system_bridge_s0_readdatavalid
	wire   [3:0] mm_interconnect_0_out_system_bridge_s0_byteenable;                          // mm_interconnect_0:out_system_bridge_s0_byteenable -> out_system_bridge:s0_byteenable
	wire  [31:0] mm_interconnect_0_button_pio_s1_writedata;                                  // mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	wire   [1:0] mm_interconnect_0_button_pio_s1_address;                                    // mm_interconnect_0:button_pio_s1_address -> button_pio:address
	wire         mm_interconnect_0_button_pio_s1_chipselect;                                 // mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	wire         mm_interconnect_0_button_pio_s1_write;                                      // mm_interconnect_0:button_pio_s1_write -> button_pio:write_n
	wire  [31:0] mm_interconnect_0_button_pio_s1_readdata;                                   // button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	wire         irq_mapper_receiver0_irq;                                                   // timer:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                   // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                   // button_pio:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                   // cpu_irq_0:ins_irq0_irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                   // fprint_irq_0:irq_out -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                   // dma_0_irq:sender0_irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                                   // dma_0_irq:sender1_irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver8_irq;                                                   // dma_0_irq:sender2_irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                                                   // dma_0_irq:sender3_irq -> irq_mapper:receiver9_irq
	wire  [31:0] cpum_d_irq_irq;                                                             // irq_mapper:sender_irq -> cpuM:d_irq
	wire         rst_controller_reset_out_reset;                                             // rst_controller:reset_out -> [button_pio:reset_n, cpuM:reset_n, cpu_irq_0:reset, dma_0_irq:reset, fprint_irq_0:reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:cpuM_reset_n_reset_bridge_in_reset_reset, out_system_bridge:reset, rst_translator:in_reset, scratchpad:reset, timer:reset_n, timestamp:reset_n]
	wire         rst_controller_reset_out_reset_req;                                         // rst_controller:reset_req -> [cpuM:reset_req, rst_translator:reset_req_in, scratchpad:reset_req]

	nios_fprint_processorM_0_cpuM cpum (
		.clk                                   (philosopher_clk_in_clk),                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                      //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                             (cpum_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpum_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpum_data_master_read),                                //                          .read
		.d_readdata                            (cpum_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpum_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpum_data_master_write),                               //                          .write
		.d_writedata                           (cpum_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpum_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpum_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpum_instruction_master_read),                         //                          .read
		.i_readdata                            (cpum_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpum_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpum_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpum_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpum_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpum_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpum_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpum_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpum_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpum_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpum_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpum_jtag_debug_module_writedata),   //                          .writedata
		.A_ci_multi_done                       (cpum_custom_instruction_master_done),                  // custom_instruction_master.done
		.A_ci_multi_result                     (cpum_custom_instruction_master_multi_result),          //                          .multi_result
		.A_ci_multi_a                          (cpum_custom_instruction_master_multi_a),               //                          .multi_a
		.A_ci_multi_b                          (cpum_custom_instruction_master_multi_b),               //                          .multi_b
		.A_ci_multi_c                          (cpum_custom_instruction_master_multi_c),               //                          .multi_c
		.A_ci_multi_clk_en                     (cpum_custom_instruction_master_clk_en),                //                          .clk_en
		.A_ci_multi_clock                      (cpum_custom_instruction_master_clk),                   //                          .clk
		.A_ci_multi_reset                      (cpum_custom_instruction_master_reset),                 //                          .reset
		.A_ci_multi_reset_req                  (cpum_custom_instruction_master_reset_req),             //                          .reset_req
		.A_ci_multi_dataa                      (cpum_custom_instruction_master_multi_dataa),           //                          .multi_dataa
		.A_ci_multi_datab                      (cpum_custom_instruction_master_multi_datab),           //                          .multi_datab
		.A_ci_multi_n                          (cpum_custom_instruction_master_multi_n),               //                          .multi_n
		.A_ci_multi_readra                     (cpum_custom_instruction_master_multi_readra),          //                          .multi_readra
		.A_ci_multi_readrb                     (cpum_custom_instruction_master_multi_readrb),          //                          .multi_readrb
		.A_ci_multi_start                      (cpum_custom_instruction_master_start),                 //                          .start
		.A_ci_multi_writerc                    (cpum_custom_instruction_master_multi_writerc),         //                          .multi_writerc
		.E_ci_combo_result                     (cpum_custom_instruction_master_result),                //                          .result
		.E_ci_combo_a                          (cpum_custom_instruction_master_a),                     //                          .a
		.E_ci_combo_b                          (cpum_custom_instruction_master_b),                     //                          .b
		.E_ci_combo_c                          (cpum_custom_instruction_master_c),                     //                          .c
		.E_ci_combo_dataa                      (cpum_custom_instruction_master_dataa),                 //                          .dataa
		.E_ci_combo_datab                      (cpum_custom_instruction_master_datab),                 //                          .datab
		.E_ci_combo_n                          (cpum_custom_instruction_master_n),                     //                          .n
		.E_ci_combo_readra                     (cpum_custom_instruction_master_readra),                //                          .readra
		.E_ci_combo_readrb                     (cpum_custom_instruction_master_readrb),                //                          .readrb
		.E_ci_combo_writerc                    (cpum_custom_instruction_master_writerc)                //                          .writerc
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (27),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) out_system_bridge (
		.clk              (philosopher_clk_in_clk),                               //   clk.clk
		.reset            (rst_controller_reset_out_reset),                       // reset.reset
		.s0_waitrequest   (mm_interconnect_0_out_system_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_out_system_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_out_system_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_out_system_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_out_system_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_out_system_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_out_system_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_out_system_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_out_system_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_out_system_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (outgoing_master_waitrequest),                          //    m0.waitrequest
		.m0_readdata      (outgoing_master_readdata),                             //      .readdata
		.m0_readdatavalid (outgoing_master_readdatavalid),                        //      .readdatavalid
		.m0_burstcount    (outgoing_master_burstcount),                           //      .burstcount
		.m0_writedata     (outgoing_master_writedata),                            //      .writedata
		.m0_address       (outgoing_master_address),                              //      .address
		.m0_write         (outgoing_master_write),                                //      .write
		.m0_read          (outgoing_master_read),                                 //      .read
		.m0_byteenable    (outgoing_master_byteenable),                           //      .byteenable
		.m0_debugaccess   (outgoing_master_debugaccess)                           //      .debugaccess
	);

	nios_fprint_processor1_0_timer timer (
		.clk        (philosopher_clk_in_clk),                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)               //   irq.irq
	);

	nios_fprint_processor1_0_jtag_uart jtag_uart (
		.clk            (philosopher_clk_in_clk),                                    //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	nios_fprint_processor1_0_button_pio button_pio (
		.clk        (philosopher_clk_in_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_button_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button_pio_s1_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                    //                 irq.irq
	);

	cpu_irq cpu_irq_0 (
		.avs_s0_address   (cpu_irq_0_s0_address),           //    s0.address
		.avs_s0_write     (cpu_irq_0_s0_write),             //      .write
		.avs_s0_writedata (cpu_irq_0_s0_writedata),         //      .writedata
		.clk              (philosopher_clk_in_clk),         // clock.clk
		.reset            (rst_controller_reset_out_reset), // reset.reset
		.ins_irq0_irq     (irq_mapper_receiver3_irq)        //  irq0.irq
	);

	nios_fprint_processor1_0_timestamp timestamp (
		.clk        (philosopher_clk_in_clk),                    //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_timestamp_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timestamp_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timestamp_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timestamp_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timestamp_s1_write),     //      .write_n
		.irq        ()                                           //   irq.irq
	);

	fprint_irq fprint_irq_0 (
		.irq_out (irq_mapper_receiver4_irq),       // interrupt_sender.irq
		.irq     (fprint_irq_0_irq_export),        //              irq.export
		.clk     (philosopher_clk_in_clk),         //            clock.clk
		.reset   (rst_controller_reset_out_reset)  //            reset.reset
	);

	altera_irq_bridge #(
		.IRQ_WIDTH (4)
	) dma_0_irq (
		.clk          (philosopher_clk_in_clk),         //          clk.clk
		.receiver_irq (dma_0_irq_receiver_irq_irq),     // receiver_irq.irq
		.reset        (rst_controller_reset_out_reset), //    clk_reset.reset
		.sender0_irq  (irq_mapper_receiver5_irq),       //  sender0_irq.irq
		.sender1_irq  (irq_mapper_receiver6_irq),       //  sender1_irq.irq
		.sender2_irq  (irq_mapper_receiver8_irq),       //  sender2_irq.irq
		.sender3_irq  (irq_mapper_receiver9_irq),       //  sender3_irq.irq
		.sender4_irq  (),                               //  (terminated)
		.sender5_irq  (),                               //  (terminated)
		.sender6_irq  (),                               //  (terminated)
		.sender7_irq  (),                               //  (terminated)
		.sender8_irq  (),                               //  (terminated)
		.sender9_irq  (),                               //  (terminated)
		.sender10_irq (),                               //  (terminated)
		.sender11_irq (),                               //  (terminated)
		.sender12_irq (),                               //  (terminated)
		.sender13_irq (),                               //  (terminated)
		.sender14_irq (),                               //  (terminated)
		.sender15_irq (),                               //  (terminated)
		.sender16_irq (),                               //  (terminated)
		.sender17_irq (),                               //  (terminated)
		.sender18_irq (),                               //  (terminated)
		.sender19_irq (),                               //  (terminated)
		.sender20_irq (),                               //  (terminated)
		.sender21_irq (),                               //  (terminated)
		.sender22_irq (),                               //  (terminated)
		.sender23_irq (),                               //  (terminated)
		.sender24_irq (),                               //  (terminated)
		.sender25_irq (),                               //  (terminated)
		.sender26_irq (),                               //  (terminated)
		.sender27_irq (),                               //  (terminated)
		.sender28_irq (),                               //  (terminated)
		.sender29_irq (),                               //  (terminated)
		.sender30_irq (),                               //  (terminated)
		.sender31_irq ()                                //  (terminated)
	);

	nios_fprint_processorM_0_scratchpad scratchpad (
		.clk        (philosopher_clk_in_clk),                     //   clk1.clk
		.address    (mm_interconnect_0_scratchpad_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_scratchpad_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_scratchpad_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_scratchpad_s1_write),      //       .write
		.readdata   (mm_interconnect_0_scratchpad_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_scratchpad_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_scratchpad_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)          //       .reset_req
	);

	nios_fprint_processor1_0_nios_custom_instr_floating_point_2_0 nios_custom_instr_floating_point_2_0 (
		.s1_dataa     (cpum_custom_instruction_master_comb_slave_translator0_ci_master_dataa),      // s1.dataa
		.s1_datab     (cpum_custom_instruction_master_comb_slave_translator0_ci_master_datab),      //   .datab
		.s1_n         (cpum_custom_instruction_master_comb_slave_translator0_ci_master_n),          //   .n
		.s1_result    (cpum_custom_instruction_master_comb_slave_translator0_ci_master_result),     //   .result
		.s2_clk       (cpum_custom_instruction_master_multi_slave_translator0_ci_master_clk),       // s2.clk
		.s2_clk_en    (cpum_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //   .clk_en
		.s2_dataa     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     //   .dataa
		.s2_datab     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //   .datab
		.s2_n         (cpum_custom_instruction_master_multi_slave_translator0_ci_master_n),         //   .n
		.s2_reset     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //   .reset
		.s2_reset_req (cpum_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //   .reset_req
		.s2_start     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_start),     //   .start
		.s2_done      (cpum_custom_instruction_master_multi_slave_translator0_ci_master_done),      //   .done
		.s2_result    (cpum_custom_instruction_master_multi_slave_translator0_ci_master_result)     //   .result
	);

	altera_customins_master_translator #(
		.SHARED_COMB_AND_MULTI (0)
	) cpum_custom_instruction_master_translator (
		.ci_slave_dataa            (cpum_custom_instruction_master_dataa),                                //        ci_slave.dataa
		.ci_slave_datab            (cpum_custom_instruction_master_datab),                                //                .datab
		.ci_slave_result           (cpum_custom_instruction_master_result),                               //                .result
		.ci_slave_n                (cpum_custom_instruction_master_n),                                    //                .n
		.ci_slave_readra           (cpum_custom_instruction_master_readra),                               //                .readra
		.ci_slave_readrb           (cpum_custom_instruction_master_readrb),                               //                .readrb
		.ci_slave_writerc          (cpum_custom_instruction_master_writerc),                              //                .writerc
		.ci_slave_a                (cpum_custom_instruction_master_a),                                    //                .a
		.ci_slave_b                (cpum_custom_instruction_master_b),                                    //                .b
		.ci_slave_c                (cpum_custom_instruction_master_c),                                    //                .c
		.ci_slave_ipending         (),                                                                    //                .ipending
		.ci_slave_estatus          (),                                                                    //                .estatus
		.ci_slave_multi_clk        (cpum_custom_instruction_master_clk),                                  //                .clk
		.ci_slave_multi_reset      (cpum_custom_instruction_master_reset),                                //                .reset
		.ci_slave_multi_clken      (cpum_custom_instruction_master_clk_en),                               //                .clk_en
		.ci_slave_multi_reset_req  (cpum_custom_instruction_master_reset_req),                            //                .reset_req
		.ci_slave_multi_start      (cpum_custom_instruction_master_start),                                //                .start
		.ci_slave_multi_done       (cpum_custom_instruction_master_done),                                 //                .done
		.ci_slave_multi_dataa      (cpum_custom_instruction_master_multi_dataa),                          //                .multi_dataa
		.ci_slave_multi_datab      (cpum_custom_instruction_master_multi_datab),                          //                .multi_datab
		.ci_slave_multi_result     (cpum_custom_instruction_master_multi_result),                         //                .multi_result
		.ci_slave_multi_n          (cpum_custom_instruction_master_multi_n),                              //                .multi_n
		.ci_slave_multi_readra     (cpum_custom_instruction_master_multi_readra),                         //                .multi_readra
		.ci_slave_multi_readrb     (cpum_custom_instruction_master_multi_readrb),                         //                .multi_readrb
		.ci_slave_multi_writerc    (cpum_custom_instruction_master_multi_writerc),                        //                .multi_writerc
		.ci_slave_multi_a          (cpum_custom_instruction_master_multi_a),                              //                .multi_a
		.ci_slave_multi_b          (cpum_custom_instruction_master_multi_b),                              //                .multi_b
		.ci_slave_multi_c          (cpum_custom_instruction_master_multi_c),                              //                .multi_c
		.comb_ci_master_dataa      (cpum_custom_instruction_master_translator_comb_ci_master_dataa),      //  comb_ci_master.dataa
		.comb_ci_master_datab      (cpum_custom_instruction_master_translator_comb_ci_master_datab),      //                .datab
		.comb_ci_master_result     (cpum_custom_instruction_master_translator_comb_ci_master_result),     //                .result
		.comb_ci_master_n          (cpum_custom_instruction_master_translator_comb_ci_master_n),          //                .n
		.comb_ci_master_readra     (cpum_custom_instruction_master_translator_comb_ci_master_readra),     //                .readra
		.comb_ci_master_readrb     (cpum_custom_instruction_master_translator_comb_ci_master_readrb),     //                .readrb
		.comb_ci_master_writerc    (cpum_custom_instruction_master_translator_comb_ci_master_writerc),    //                .writerc
		.comb_ci_master_a          (cpum_custom_instruction_master_translator_comb_ci_master_a),          //                .a
		.comb_ci_master_b          (cpum_custom_instruction_master_translator_comb_ci_master_b),          //                .b
		.comb_ci_master_c          (cpum_custom_instruction_master_translator_comb_ci_master_c),          //                .c
		.comb_ci_master_ipending   (cpum_custom_instruction_master_translator_comb_ci_master_ipending),   //                .ipending
		.comb_ci_master_estatus    (cpum_custom_instruction_master_translator_comb_ci_master_estatus),    //                .estatus
		.multi_ci_master_clk       (cpum_custom_instruction_master_translator_multi_ci_master_clk),       // multi_ci_master.clk
		.multi_ci_master_reset     (cpum_custom_instruction_master_translator_multi_ci_master_reset),     //                .reset
		.multi_ci_master_clken     (cpum_custom_instruction_master_translator_multi_ci_master_clk_en),    //                .clk_en
		.multi_ci_master_reset_req (cpum_custom_instruction_master_translator_multi_ci_master_reset_req), //                .reset_req
		.multi_ci_master_start     (cpum_custom_instruction_master_translator_multi_ci_master_start),     //                .start
		.multi_ci_master_done      (cpum_custom_instruction_master_translator_multi_ci_master_done),      //                .done
		.multi_ci_master_dataa     (cpum_custom_instruction_master_translator_multi_ci_master_dataa),     //                .dataa
		.multi_ci_master_datab     (cpum_custom_instruction_master_translator_multi_ci_master_datab),     //                .datab
		.multi_ci_master_result    (cpum_custom_instruction_master_translator_multi_ci_master_result),    //                .result
		.multi_ci_master_n         (cpum_custom_instruction_master_translator_multi_ci_master_n),         //                .n
		.multi_ci_master_readra    (cpum_custom_instruction_master_translator_multi_ci_master_readra),    //                .readra
		.multi_ci_master_readrb    (cpum_custom_instruction_master_translator_multi_ci_master_readrb),    //                .readrb
		.multi_ci_master_writerc   (cpum_custom_instruction_master_translator_multi_ci_master_writerc),   //                .writerc
		.multi_ci_master_a         (cpum_custom_instruction_master_translator_multi_ci_master_a),         //                .a
		.multi_ci_master_b         (cpum_custom_instruction_master_translator_multi_ci_master_b),         //                .b
		.multi_ci_master_c         (cpum_custom_instruction_master_translator_multi_ci_master_c)          //                .c
	);

	nios_fprint_processor1_0_cpu1_custom_instruction_master_comb_xconnect cpum_custom_instruction_master_comb_xconnect (
		.ci_slave_dataa      (cpum_custom_instruction_master_translator_comb_ci_master_dataa),    //   ci_slave.dataa
		.ci_slave_datab      (cpum_custom_instruction_master_translator_comb_ci_master_datab),    //           .datab
		.ci_slave_result     (cpum_custom_instruction_master_translator_comb_ci_master_result),   //           .result
		.ci_slave_n          (cpum_custom_instruction_master_translator_comb_ci_master_n),        //           .n
		.ci_slave_readra     (cpum_custom_instruction_master_translator_comb_ci_master_readra),   //           .readra
		.ci_slave_readrb     (cpum_custom_instruction_master_translator_comb_ci_master_readrb),   //           .readrb
		.ci_slave_writerc    (cpum_custom_instruction_master_translator_comb_ci_master_writerc),  //           .writerc
		.ci_slave_a          (cpum_custom_instruction_master_translator_comb_ci_master_a),        //           .a
		.ci_slave_b          (cpum_custom_instruction_master_translator_comb_ci_master_b),        //           .b
		.ci_slave_c          (cpum_custom_instruction_master_translator_comb_ci_master_c),        //           .c
		.ci_slave_ipending   (cpum_custom_instruction_master_translator_comb_ci_master_ipending), //           .ipending
		.ci_slave_estatus    (cpum_custom_instruction_master_translator_comb_ci_master_estatus),  //           .estatus
		.ci_master0_dataa    (cpum_custom_instruction_master_comb_xconnect_ci_master0_dataa),     // ci_master0.dataa
		.ci_master0_datab    (cpum_custom_instruction_master_comb_xconnect_ci_master0_datab),     //           .datab
		.ci_master0_result   (cpum_custom_instruction_master_comb_xconnect_ci_master0_result),    //           .result
		.ci_master0_n        (cpum_custom_instruction_master_comb_xconnect_ci_master0_n),         //           .n
		.ci_master0_readra   (cpum_custom_instruction_master_comb_xconnect_ci_master0_readra),    //           .readra
		.ci_master0_readrb   (cpum_custom_instruction_master_comb_xconnect_ci_master0_readrb),    //           .readrb
		.ci_master0_writerc  (cpum_custom_instruction_master_comb_xconnect_ci_master0_writerc),   //           .writerc
		.ci_master0_a        (cpum_custom_instruction_master_comb_xconnect_ci_master0_a),         //           .a
		.ci_master0_b        (cpum_custom_instruction_master_comb_xconnect_ci_master0_b),         //           .b
		.ci_master0_c        (cpum_custom_instruction_master_comb_xconnect_ci_master0_c),         //           .c
		.ci_master0_ipending (cpum_custom_instruction_master_comb_xconnect_ci_master0_ipending),  //           .ipending
		.ci_master0_estatus  (cpum_custom_instruction_master_comb_xconnect_ci_master0_estatus)    //           .estatus
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (4),
		.USE_DONE         (0),
		.NUM_FIXED_CYCLES (0)
	) cpum_custom_instruction_master_comb_slave_translator0 (
		.ci_slave_dataa      (cpum_custom_instruction_master_comb_xconnect_ci_master0_dataa),          //  ci_slave.dataa
		.ci_slave_datab      (cpum_custom_instruction_master_comb_xconnect_ci_master0_datab),          //          .datab
		.ci_slave_result     (cpum_custom_instruction_master_comb_xconnect_ci_master0_result),         //          .result
		.ci_slave_n          (cpum_custom_instruction_master_comb_xconnect_ci_master0_n),              //          .n
		.ci_slave_readra     (cpum_custom_instruction_master_comb_xconnect_ci_master0_readra),         //          .readra
		.ci_slave_readrb     (cpum_custom_instruction_master_comb_xconnect_ci_master0_readrb),         //          .readrb
		.ci_slave_writerc    (cpum_custom_instruction_master_comb_xconnect_ci_master0_writerc),        //          .writerc
		.ci_slave_a          (cpum_custom_instruction_master_comb_xconnect_ci_master0_a),              //          .a
		.ci_slave_b          (cpum_custom_instruction_master_comb_xconnect_ci_master0_b),              //          .b
		.ci_slave_c          (cpum_custom_instruction_master_comb_xconnect_ci_master0_c),              //          .c
		.ci_slave_ipending   (cpum_custom_instruction_master_comb_xconnect_ci_master0_ipending),       //          .ipending
		.ci_slave_estatus    (cpum_custom_instruction_master_comb_xconnect_ci_master0_estatus),        //          .estatus
		.ci_master_dataa     (cpum_custom_instruction_master_comb_slave_translator0_ci_master_dataa),  // ci_master.dataa
		.ci_master_datab     (cpum_custom_instruction_master_comb_slave_translator0_ci_master_datab),  //          .datab
		.ci_master_result    (cpum_custom_instruction_master_comb_slave_translator0_ci_master_result), //          .result
		.ci_master_n         (cpum_custom_instruction_master_comb_slave_translator0_ci_master_n),      //          .n
		.ci_master_readra    (),                                                                       // (terminated)
		.ci_master_readrb    (),                                                                       // (terminated)
		.ci_master_writerc   (),                                                                       // (terminated)
		.ci_master_a         (),                                                                       // (terminated)
		.ci_master_b         (),                                                                       // (terminated)
		.ci_master_c         (),                                                                       // (terminated)
		.ci_master_ipending  (),                                                                       // (terminated)
		.ci_master_estatus   (),                                                                       // (terminated)
		.ci_master_clk       (),                                                                       // (terminated)
		.ci_master_clken     (),                                                                       // (terminated)
		.ci_master_reset_req (),                                                                       // (terminated)
		.ci_master_reset     (),                                                                       // (terminated)
		.ci_master_start     (),                                                                       // (terminated)
		.ci_master_done      (1'b0),                                                                   // (terminated)
		.ci_slave_clk        (1'b0),                                                                   // (terminated)
		.ci_slave_clken      (1'b0),                                                                   // (terminated)
		.ci_slave_reset_req  (1'b0),                                                                   // (terminated)
		.ci_slave_reset      (1'b0),                                                                   // (terminated)
		.ci_slave_start      (1'b0),                                                                   // (terminated)
		.ci_slave_done       ()                                                                        // (terminated)
	);

	nios_fprint_processor1_0_cpu1_custom_instruction_master_multi_xconnect cpum_custom_instruction_master_multi_xconnect (
		.ci_slave_dataa       (cpum_custom_instruction_master_translator_multi_ci_master_dataa),     //   ci_slave.dataa
		.ci_slave_datab       (cpum_custom_instruction_master_translator_multi_ci_master_datab),     //           .datab
		.ci_slave_result      (cpum_custom_instruction_master_translator_multi_ci_master_result),    //           .result
		.ci_slave_n           (cpum_custom_instruction_master_translator_multi_ci_master_n),         //           .n
		.ci_slave_readra      (cpum_custom_instruction_master_translator_multi_ci_master_readra),    //           .readra
		.ci_slave_readrb      (cpum_custom_instruction_master_translator_multi_ci_master_readrb),    //           .readrb
		.ci_slave_writerc     (cpum_custom_instruction_master_translator_multi_ci_master_writerc),   //           .writerc
		.ci_slave_a           (cpum_custom_instruction_master_translator_multi_ci_master_a),         //           .a
		.ci_slave_b           (cpum_custom_instruction_master_translator_multi_ci_master_b),         //           .b
		.ci_slave_c           (cpum_custom_instruction_master_translator_multi_ci_master_c),         //           .c
		.ci_slave_ipending    (),                                                                    //           .ipending
		.ci_slave_estatus     (),                                                                    //           .estatus
		.ci_slave_clk         (cpum_custom_instruction_master_translator_multi_ci_master_clk),       //           .clk
		.ci_slave_reset       (cpum_custom_instruction_master_translator_multi_ci_master_reset),     //           .reset
		.ci_slave_clken       (cpum_custom_instruction_master_translator_multi_ci_master_clk_en),    //           .clk_en
		.ci_slave_reset_req   (cpum_custom_instruction_master_translator_multi_ci_master_reset_req), //           .reset_req
		.ci_slave_start       (cpum_custom_instruction_master_translator_multi_ci_master_start),     //           .start
		.ci_slave_done        (cpum_custom_instruction_master_translator_multi_ci_master_done),      //           .done
		.ci_master0_dataa     (cpum_custom_instruction_master_multi_xconnect_ci_master0_dataa),      // ci_master0.dataa
		.ci_master0_datab     (cpum_custom_instruction_master_multi_xconnect_ci_master0_datab),      //           .datab
		.ci_master0_result    (cpum_custom_instruction_master_multi_xconnect_ci_master0_result),     //           .result
		.ci_master0_n         (cpum_custom_instruction_master_multi_xconnect_ci_master0_n),          //           .n
		.ci_master0_readra    (cpum_custom_instruction_master_multi_xconnect_ci_master0_readra),     //           .readra
		.ci_master0_readrb    (cpum_custom_instruction_master_multi_xconnect_ci_master0_readrb),     //           .readrb
		.ci_master0_writerc   (cpum_custom_instruction_master_multi_xconnect_ci_master0_writerc),    //           .writerc
		.ci_master0_a         (cpum_custom_instruction_master_multi_xconnect_ci_master0_a),          //           .a
		.ci_master0_b         (cpum_custom_instruction_master_multi_xconnect_ci_master0_b),          //           .b
		.ci_master0_c         (cpum_custom_instruction_master_multi_xconnect_ci_master0_c),          //           .c
		.ci_master0_ipending  (cpum_custom_instruction_master_multi_xconnect_ci_master0_ipending),   //           .ipending
		.ci_master0_estatus   (cpum_custom_instruction_master_multi_xconnect_ci_master0_estatus),    //           .estatus
		.ci_master0_clk       (cpum_custom_instruction_master_multi_xconnect_ci_master0_clk),        //           .clk
		.ci_master0_reset     (cpum_custom_instruction_master_multi_xconnect_ci_master0_reset),      //           .reset
		.ci_master0_clken     (cpum_custom_instruction_master_multi_xconnect_ci_master0_clk_en),     //           .clk_en
		.ci_master0_reset_req (cpum_custom_instruction_master_multi_xconnect_ci_master0_reset_req),  //           .reset_req
		.ci_master0_start     (cpum_custom_instruction_master_multi_xconnect_ci_master0_start),      //           .start
		.ci_master0_done      (cpum_custom_instruction_master_multi_xconnect_ci_master0_done)        //           .done
	);

	altera_customins_slave_translator #(
		.N_WIDTH          (3),
		.USE_DONE         (1),
		.NUM_FIXED_CYCLES (1)
	) cpum_custom_instruction_master_multi_slave_translator0 (
		.ci_slave_dataa      (cpum_custom_instruction_master_multi_xconnect_ci_master0_dataa),             //  ci_slave.dataa
		.ci_slave_datab      (cpum_custom_instruction_master_multi_xconnect_ci_master0_datab),             //          .datab
		.ci_slave_result     (cpum_custom_instruction_master_multi_xconnect_ci_master0_result),            //          .result
		.ci_slave_n          (cpum_custom_instruction_master_multi_xconnect_ci_master0_n),                 //          .n
		.ci_slave_readra     (cpum_custom_instruction_master_multi_xconnect_ci_master0_readra),            //          .readra
		.ci_slave_readrb     (cpum_custom_instruction_master_multi_xconnect_ci_master0_readrb),            //          .readrb
		.ci_slave_writerc    (cpum_custom_instruction_master_multi_xconnect_ci_master0_writerc),           //          .writerc
		.ci_slave_a          (cpum_custom_instruction_master_multi_xconnect_ci_master0_a),                 //          .a
		.ci_slave_b          (cpum_custom_instruction_master_multi_xconnect_ci_master0_b),                 //          .b
		.ci_slave_c          (cpum_custom_instruction_master_multi_xconnect_ci_master0_c),                 //          .c
		.ci_slave_ipending   (cpum_custom_instruction_master_multi_xconnect_ci_master0_ipending),          //          .ipending
		.ci_slave_estatus    (cpum_custom_instruction_master_multi_xconnect_ci_master0_estatus),           //          .estatus
		.ci_slave_clk        (cpum_custom_instruction_master_multi_xconnect_ci_master0_clk),               //          .clk
		.ci_slave_clken      (cpum_custom_instruction_master_multi_xconnect_ci_master0_clk_en),            //          .clk_en
		.ci_slave_reset_req  (cpum_custom_instruction_master_multi_xconnect_ci_master0_reset_req),         //          .reset_req
		.ci_slave_reset      (cpum_custom_instruction_master_multi_xconnect_ci_master0_reset),             //          .reset
		.ci_slave_start      (cpum_custom_instruction_master_multi_xconnect_ci_master0_start),             //          .start
		.ci_slave_done       (cpum_custom_instruction_master_multi_xconnect_ci_master0_done),              //          .done
		.ci_master_dataa     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_dataa),     // ci_master.dataa
		.ci_master_datab     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_datab),     //          .datab
		.ci_master_result    (cpum_custom_instruction_master_multi_slave_translator0_ci_master_result),    //          .result
		.ci_master_n         (cpum_custom_instruction_master_multi_slave_translator0_ci_master_n),         //          .n
		.ci_master_clk       (cpum_custom_instruction_master_multi_slave_translator0_ci_master_clk),       //          .clk
		.ci_master_clken     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_clk_en),    //          .clk_en
		.ci_master_reset_req (cpum_custom_instruction_master_multi_slave_translator0_ci_master_reset_req), //          .reset_req
		.ci_master_reset     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_reset),     //          .reset
		.ci_master_start     (cpum_custom_instruction_master_multi_slave_translator0_ci_master_start),     //          .start
		.ci_master_done      (cpum_custom_instruction_master_multi_slave_translator0_ci_master_done),      //          .done
		.ci_master_readra    (),                                                                           // (terminated)
		.ci_master_readrb    (),                                                                           // (terminated)
		.ci_master_writerc   (),                                                                           // (terminated)
		.ci_master_a         (),                                                                           // (terminated)
		.ci_master_b         (),                                                                           // (terminated)
		.ci_master_c         (),                                                                           // (terminated)
		.ci_master_ipending  (),                                                                           // (terminated)
		.ci_master_estatus   ()                                                                            // (terminated)
	);

	nios_fprint_processorM_0_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                              (philosopher_clk_in_clk),                                    //                            clk_clk.clk
		.cpuM_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // cpuM_reset_n_reset_bridge_in_reset.reset
		.cpuM_data_master_address                 (cpum_data_master_address),                                  //                   cpuM_data_master.address
		.cpuM_data_master_waitrequest             (cpum_data_master_waitrequest),                              //                                   .waitrequest
		.cpuM_data_master_byteenable              (cpum_data_master_byteenable),                               //                                   .byteenable
		.cpuM_data_master_read                    (cpum_data_master_read),                                     //                                   .read
		.cpuM_data_master_readdata                (cpum_data_master_readdata),                                 //                                   .readdata
		.cpuM_data_master_write                   (cpum_data_master_write),                                    //                                   .write
		.cpuM_data_master_writedata               (cpum_data_master_writedata),                                //                                   .writedata
		.cpuM_data_master_debugaccess             (cpum_data_master_debugaccess),                              //                                   .debugaccess
		.cpuM_instruction_master_address          (cpum_instruction_master_address),                           //            cpuM_instruction_master.address
		.cpuM_instruction_master_waitrequest      (cpum_instruction_master_waitrequest),                       //                                   .waitrequest
		.cpuM_instruction_master_read             (cpum_instruction_master_read),                              //                                   .read
		.cpuM_instruction_master_readdata         (cpum_instruction_master_readdata),                          //                                   .readdata
		.cpuM_instruction_master_readdatavalid    (cpum_instruction_master_readdatavalid),                     //                                   .readdatavalid
		.button_pio_s1_address                    (mm_interconnect_0_button_pio_s1_address),                   //                      button_pio_s1.address
		.button_pio_s1_write                      (mm_interconnect_0_button_pio_s1_write),                     //                                   .write
		.button_pio_s1_readdata                   (mm_interconnect_0_button_pio_s1_readdata),                  //                                   .readdata
		.button_pio_s1_writedata                  (mm_interconnect_0_button_pio_s1_writedata),                 //                                   .writedata
		.button_pio_s1_chipselect                 (mm_interconnect_0_button_pio_s1_chipselect),                //                                   .chipselect
		.cpuM_jtag_debug_module_address           (mm_interconnect_0_cpum_jtag_debug_module_address),          //             cpuM_jtag_debug_module.address
		.cpuM_jtag_debug_module_write             (mm_interconnect_0_cpum_jtag_debug_module_write),            //                                   .write
		.cpuM_jtag_debug_module_read              (mm_interconnect_0_cpum_jtag_debug_module_read),             //                                   .read
		.cpuM_jtag_debug_module_readdata          (mm_interconnect_0_cpum_jtag_debug_module_readdata),         //                                   .readdata
		.cpuM_jtag_debug_module_writedata         (mm_interconnect_0_cpum_jtag_debug_module_writedata),        //                                   .writedata
		.cpuM_jtag_debug_module_byteenable        (mm_interconnect_0_cpum_jtag_debug_module_byteenable),       //                                   .byteenable
		.cpuM_jtag_debug_module_waitrequest       (mm_interconnect_0_cpum_jtag_debug_module_waitrequest),      //                                   .waitrequest
		.cpuM_jtag_debug_module_debugaccess       (mm_interconnect_0_cpum_jtag_debug_module_debugaccess),      //                                   .debugaccess
		.jtag_uart_avalon_jtag_slave_address      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                   .write
		.jtag_uart_avalon_jtag_slave_read         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                   .read
		.jtag_uart_avalon_jtag_slave_readdata     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                   .chipselect
		.out_system_bridge_s0_address             (mm_interconnect_0_out_system_bridge_s0_address),            //               out_system_bridge_s0.address
		.out_system_bridge_s0_write               (mm_interconnect_0_out_system_bridge_s0_write),              //                                   .write
		.out_system_bridge_s0_read                (mm_interconnect_0_out_system_bridge_s0_read),               //                                   .read
		.out_system_bridge_s0_readdata            (mm_interconnect_0_out_system_bridge_s0_readdata),           //                                   .readdata
		.out_system_bridge_s0_writedata           (mm_interconnect_0_out_system_bridge_s0_writedata),          //                                   .writedata
		.out_system_bridge_s0_burstcount          (mm_interconnect_0_out_system_bridge_s0_burstcount),         //                                   .burstcount
		.out_system_bridge_s0_byteenable          (mm_interconnect_0_out_system_bridge_s0_byteenable),         //                                   .byteenable
		.out_system_bridge_s0_readdatavalid       (mm_interconnect_0_out_system_bridge_s0_readdatavalid),      //                                   .readdatavalid
		.out_system_bridge_s0_waitrequest         (mm_interconnect_0_out_system_bridge_s0_waitrequest),        //                                   .waitrequest
		.out_system_bridge_s0_debugaccess         (mm_interconnect_0_out_system_bridge_s0_debugaccess),        //                                   .debugaccess
		.scratchpad_s1_address                    (mm_interconnect_0_scratchpad_s1_address),                   //                      scratchpad_s1.address
		.scratchpad_s1_write                      (mm_interconnect_0_scratchpad_s1_write),                     //                                   .write
		.scratchpad_s1_readdata                   (mm_interconnect_0_scratchpad_s1_readdata),                  //                                   .readdata
		.scratchpad_s1_writedata                  (mm_interconnect_0_scratchpad_s1_writedata),                 //                                   .writedata
		.scratchpad_s1_byteenable                 (mm_interconnect_0_scratchpad_s1_byteenable),                //                                   .byteenable
		.scratchpad_s1_chipselect                 (mm_interconnect_0_scratchpad_s1_chipselect),                //                                   .chipselect
		.scratchpad_s1_clken                      (mm_interconnect_0_scratchpad_s1_clken),                     //                                   .clken
		.timer_s1_address                         (mm_interconnect_0_timer_s1_address),                        //                           timer_s1.address
		.timer_s1_write                           (mm_interconnect_0_timer_s1_write),                          //                                   .write
		.timer_s1_readdata                        (mm_interconnect_0_timer_s1_readdata),                       //                                   .readdata
		.timer_s1_writedata                       (mm_interconnect_0_timer_s1_writedata),                      //                                   .writedata
		.timer_s1_chipselect                      (mm_interconnect_0_timer_s1_chipselect),                     //                                   .chipselect
		.timestamp_s1_address                     (mm_interconnect_0_timestamp_s1_address),                    //                       timestamp_s1.address
		.timestamp_s1_write                       (mm_interconnect_0_timestamp_s1_write),                      //                                   .write
		.timestamp_s1_readdata                    (mm_interconnect_0_timestamp_s1_readdata),                   //                                   .readdata
		.timestamp_s1_writedata                   (mm_interconnect_0_timestamp_s1_writedata),                  //                                   .writedata
		.timestamp_s1_chipselect                  (mm_interconnect_0_timestamp_s1_chipselect)                  //                                   .chipselect
	);

	nios_fprint_processorM_0_irq_mapper irq_mapper (
		.clk           (philosopher_clk_in_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (),                               // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.receiver9_irq (irq_mapper_receiver9_irq),       // receiver9.irq
		.sender_irq    (cpum_d_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (philosopher_clk_in_clk),             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
